CircuitMaker Text
5.6
Probes: 1
U2A_1
Transient Analysis
0 316 79 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 110 10
176 83 1022 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 2 1
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 179 457 276
9961490 0
0
6 Title:
5 Name:
0
0
0
19
7 Ground~
168 96 228 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5130 0 0
2
41966 0
0
11 Signal Gen~
195 29 188 0 64 64
0 11 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1056964608 0 1094713344
0 814313567 814313567 1065353216 1073741824 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 0.5 0 12 0 1e-09 1e-09 1 2 0
0 0 0 0 0 0 0 0 0 0
0
0 0 1344 0
5 0/12V
-18 -30 17 -22
2 V1
-8 -40 6 -32
4 F/!B
-13 -44 15 -36
0
37 %D %1 %2 DC 0 PULSE(0 12 0 1n 1n 1 2)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
391 0 0
2
41966 1
0
14 Opto Isolator~
173 149 195 0 4 9
0 12 2 3 2
0
0 0 880 0
6 OP4N25
-20 20 22 28
2 U1
-6 -29 8 -21
0
0
17 %D %1 %2 %3 %4 %S
0
0
4 DIP6
9

0 1 2 5 4 1 2 5 4 0
88 0 0 0 1 0 0 0
1 U
3124 0 0
2
41966 2
0
7 Ground~
168 186 228 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3421 0 0
2
41966 3
0
8 Op-Amp5~
219 280 80 0 5 11
0 5 7 9 8 6
0
0 0 832 0
5 TL082
9 -12 44 -4
3 U2A
16 -22 37 -14
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 1 0
1 U
8157 0 0
2
41966 4
0
7 Ground~
168 251 228 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5572 0 0
2
41966 5
0
7 N-JFET~
219 243 132 0 3 7
0 5 3 2
0
0 0 832 0
6 2N4393
12 0 54 8
2 Q1
26 -10 40 -2
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-18
7

0 2 3 1 2 3 1 0
74 0 0 0 1 0 0 0
1 Q
8901 0 0
2
41966 6
0
2 +V
167 221 232 0 1 3
0 4
0
0 0 53600 180
4 -15V
-13 1 15 9
2 V2
-6 -9 8 -1
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7361 0 0
2
41966 7
0
7 Ground~
168 176 140 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4747 0 0
2
41966 8
0
11 Signal Gen~
195 29 85 0 64 64
0 10 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1073741824 0 1092616192
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 2 0 10 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
7 -10/10V
-25 -30 24 -22
2 V3
-8 -40 6 -32
0
0
36 %D %1 %2 DC 0 SIN(0 10 2 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
972 0 0
2
41966 9
0
7 Ground~
168 137 140 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3472 0 0
2
41966 10
0
2 +V
167 280 58 0 1 3
0 9
0
0 0 53600 0
4 +15V
-12 -14 16 -6
2 V4
-5 -24 9 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9998 0 0
2
41966 11
0
2 +V
167 280 109 0 1 3
0 8
0
0 0 53600 180
4 -15V
-14 0 14 8
2 V5
-7 -10 7 -2
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3536 0 0
2
41966 12
0
11 Resistor:A~
219 94 183 0 2 5
0 12 11
0
0 0 864 180
3 560
-11 -14 10 -6
2 R1
-8 -24 6 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4597 0 0
2
41966 13
0
11 Resistor:A~
219 221 157 0 3 5
0 4 3 1
0
0 0 864 90
3 20k
7 0 28 8
2 R2
10 -10 24 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3835 0 0
2
41966 14
0
11 Resistor:A~
219 176 110 0 3 5
0 2 10 -1
0
0 0 864 90
3 10k
-28 1 -7 9
2 R3
-25 -9 -11 -1
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3670 0 0
2
41966 15
0
11 Resistor:A~
219 223 86 0 2 5
0 10 5
0
0 0 864 0
3 51k
-11 18 10 26
2 R4
-8 8 6 16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5616 0 0
2
41966 16
0
11 Resistor:A~
219 223 74 0 2 5
0 10 7
0
0 0 864 0
3 51k
-10 -14 11 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9323 0 0
2
41966 17
0
11 Resistor:A~
219 280 19 0 2 5
0 7 6
0
0 0 864 0
3 51k
-12 9 9 17
2 R6
-11 -14 3 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
317 0 0
2
41966 18
0
21
1 0 2 0 0 4096 0 1 0 0 19 2
96 222
96 207
3 0 3 0 0 8320 0 3 0 0 4 4
175 183
200 183
200 132
221 132
1 1 4 0 0 4224 0 8 15 0 0 2
221 217
221 175
2 2 3 0 0 0 0 15 7 0 0 3
221 139
221 132
230 132
1 3 2 0 0 4096 0 6 7 0 0 2
251 222
251 150
0 1 5 0 0 4224 0 0 7 17 0 2
251 86
251 114
2 5 6 0 0 8320 0 19 5 0 0 4
298 19
328 19
328 80
298 80
1 0 7 0 0 8320 0 19 0 0 16 3
262 19
251 19
251 74
4 1 8 0 0 4224 0 5 13 0 0 2
280 93
280 94
3 1 9 0 0 0 0 5 12 0 0 2
280 67
280 67
1 1 2 0 0 0 0 9 16 0 0 2
176 134
176 128
2 0 10 0 0 4096 0 16 0 0 13 2
176 92
176 80
1 0 10 0 0 4224 0 10 0 0 14 2
60 80
197 80
1 1 10 0 0 0 0 17 18 0 0 4
205 86
197 86
197 74
205 74
1 2 2 0 0 8320 0 11 10 0 0 3
137 134
137 90
60 90
2 2 7 0 0 0 0 18 5 0 0 2
241 74
262 74
2 1 5 0 0 0 0 17 5 0 0 2
241 86
262 86
1 4 2 0 0 0 0 4 3 0 0 3
186 222
186 207
175 207
2 2 2 0 0 0 0 3 2 0 0 4
121 207
71 207
71 193
60 193
1 2 11 0 0 4224 0 2 14 0 0 2
60 183
76 183
1 1 12 0 0 4224 0 14 3 0 0 2
112 183
121 183
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 10 0.02 0.02
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

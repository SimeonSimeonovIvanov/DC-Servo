CircuitMaker Text
5.6
Probes: 1
R5_2
Transient Analysis
0 406 114 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 170 10
176 79 1918 540
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 2 0
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
2 2 0.500000 0.500000
344 175 2086 645
9961490 0
0
6 Title:
5 Name:
0
0
0
17
7 Ground~
168 339 72 0 1 3
0 2
0
0 0 53360 270
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5130 0 0
2
5.89666e-315 0
0
2 +V
167 365 57 0 1 3
0 8
0
0 0 53616 0
3 15V
-10 -13 11 -5
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
391 0 0
2
5.89666e-315 5.30499e-315
0
2 +V
167 365 108 0 1 3
0 7
0
0 0 53616 180
4 -15V
-14 0 14 8
2 V3
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3124 0 0
2
5.89666e-315 5.26354e-315
0
10 Op-Amp5:A~
219 365 79 0 5 11
0 2 6 8 7 5
0
0 0 848 0
5 TL082
7 -19 42 -11
2 U2
19 -29 33 -21
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 0 0 0
1 U
3421 0 0
2
5.89666e-315 0
0
7 Ground~
168 284 121 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8157 0 0
2
5.89666e-315 0
0
10 Capacitor~
219 284 104 0 2 5
0 2 9
0
0 0 848 90
5 4.7pF
10 0 45 8
2 C1
22 -10 36 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5572 0 0
2
5.89666e-315 0
0
10 Op-Amp5:A~
219 136 169 0 5 11
0 13 4 12 11 3
0
0 0 848 0
5 TL082
7 -19 42 -11
2 U1
19 -29 33 -21
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 0 0 0
1 U
8901 0 0
2
5.89666e-315 5.37752e-315
0
2 +V
167 136 198 0 1 3
0 11
0
0 0 53616 180
4 -15V
-14 0 14 8
2 V5
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7361 0 0
2
5.89666e-315 5.36716e-315
0
7 Ground~
168 172 121 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4747 0 0
2
5.89666e-315 5.3568e-315
0
11 Signal Gen~
195 115 90 0 64 64
0 10 2 2 86 -10 10 0 0 0
0 0 0 0 0 0 0 1148846080 1075838976 1075838976
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 1000 2.5 2.5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
4 0/5V
-14 -30 14 -22
2 V2
-7 -40 7 -32
0
0
33 %D %1 %2 DC 0 SIN(2.5 2.5 1k 0 0)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
972 0 0
2
5.89666e-315 5.34643e-315
0
2 +V
167 136 147 0 1 3
0 12
0
0 0 53616 0
3 15V
-10 -13 11 -5
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3472 0 0
2
5.89666e-315 5.32571e-315
0
2 +V
167 83 165 0 1 3
0 13
0
0 0 54128 90
4 2.5V
-11 4 17 12
4 Ilim
-12 -18 16 -10
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9998 0 0
2
5.89666e-315 5.30499e-315
0
9 Schottky~
219 205 169 0 2 5
0 4 3
0
0 0 848 180
6 1N5828
-22 -18 20 -10
2 D1
-8 -28 6 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3536 0 0
2
5.89666e-315 0
0
11 Resistor:A~
219 367 152 0 2 5
0 6 5
0
0 0 880 0
2 2k
-8 -14 6 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4597 0 0
2
5.89666e-315 0
0
11 Resistor:A~
219 310 85 0 2 5
0 9 6
0
0 0 880 0
2 1k
-8 -14 6 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3835 0 0
2
5.89666e-315 0
0
11 Resistor:A~
219 198 85 0 2 5
0 10 4
0
0 0 880 0
2 1k
-8 -14 6 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3670 0 0
2
5.89666e-315 0
0
11 Resistor:A~
219 258 85 0 2 5
0 4 9
0
0 0 880 0
2 1k
-8 -14 6 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5616 0 0
2
5.89666e-315 5.38788e-315
0
18
2 5 3 0 0 4224 0 13 7 0 0 2
191 169
154 169
2 0 4 0 0 12416 0 7 0 0 12 5
118 175
108 175
108 217
229 217
229 169
1 1 2 0 0 4096 0 1 4 0 0 2
346 73
347 73
5 2 5 0 0 8320 0 4 14 0 0 4
383 79
405 79
405 152
385 152
2 0 6 0 0 4096 0 4 0 0 6 2
347 85
336 85
1 2 6 0 0 8320 0 14 15 0 0 4
349 152
336 152
336 85
328 85
4 1 7 0 0 4224 0 4 3 0 0 2
365 92
365 93
3 1 8 0 0 0 0 4 2 0 0 2
365 66
365 66
1 1 2 0 0 4096 0 5 6 0 0 2
284 115
284 113
2 0 9 0 0 4096 0 6 0 0 11 2
284 95
284 85
1 2 9 0 0 4224 0 15 17 0 0 2
292 85
276 85
1 1 4 0 0 0 0 13 17 0 0 5
214 169
229 169
229 85
228 85
240 85
1 2 2 0 0 8320 0 9 10 0 0 3
172 115
172 95
146 95
0 2 4 0 0 0 0 0 16 12 0 2
229 85
216 85
1 1 10 0 0 4224 0 10 16 0 0 2
146 85
180 85
4 1 11 0 0 4224 0 7 8 0 0 2
136 182
136 183
3 1 12 0 0 0 0 7 11 0 0 2
136 156
136 156
1 1 13 0 0 4224 0 7 12 0 0 2
118 163
94 163
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-06 2e-06
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 250 10
176 83 1022 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 2 0
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 179 457 276
42991634 0
0
6 Title:
5 Name:
0
0
0
8
13 Logic Switch~
5 92 23 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 20848 270
2 5V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5776 0 0
2
5.89683e-315 5.37752e-315
0
13 Logic Switch~
5 92 145 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 20848 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7207 0 0
2
5.89683e-315 5.36716e-315
0
13 Logic Switch~
5 14 62 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21872 0
2 5V
-6 -16 8 -8
2 V3
-6 -31 8 -23
4 A_IN
-13 -36 15 -28
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4459 0 0
2
5.89683e-315 5.3568e-315
0
13 Logic Switch~
5 14 184 0 1 11
0 2
0
0 0 21872 0
2 0V
-6 -16 8 -8
2 V4
-6 -31 8 -23
4 B_IN
-13 -36 15 -28
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3760 0 0
2
5.89683e-315 5.34643e-315
0
5 7474~
219 92 220 0 6 22
0 4 2 5 2 8 3
0
0 0 4720 0
4 7474
7 -60 35 -52
3 U2B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 4 0
1 U
754 0 0
2
5.89683e-315 5.32571e-315
0
5 7474~
219 92 98 0 6 22
0 6 5 2 5 9 7
0
0 0 4720 0
4 7474
7 -60 35 -52
3 U2A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 4 0
1 U
9767 0 0
2
5.89683e-315 5.30499e-315
0
14 Logic Display~
6 149 58 0 1 2
10 7
0
0 0 54896 270
6 100MEG
3 -16 45 -8
2 L1
-5 -15 9 -7
2 UP
-8 -35 6 -27
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7978 0 0
2
5.89683e-315 5.26354e-315
0
14 Logic Display~
6 149 180 0 1 2
10 3
0
0 0 54896 270
6 100MEG
3 -16 45 -8
2 L2
-5 -15 9 -7
4 DOWN
-15 -35 13 -27
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3142 0 0
2
5.89683e-315 0
0
10
3 0 2 0 0 8320 0 6 0 0 2 3
68 80
48 80
48 184
1 0 2 0 0 0 0 4 0 0 5 2
26 184
60 184
1 6 3 0 0 4224 0 8 5 0 0 2
133 184
116 184
1 1 4 0 0 0 0 2 5 0 0 2
92 157
92 157
4 2 2 0 0 0 0 5 5 0 0 5
92 232
92 238
60 238
60 184
68 184
4 0 5 0 0 12288 0 6 0 0 9 4
92 110
92 116
60 116
60 62
1 1 6 0 0 0 0 6 1 0 0 2
92 35
92 35
1 0 5 0 0 0 0 3 0 0 9 2
26 62
37 62
2 3 5 0 0 8320 0 6 5 0 0 4
68 62
37 62
37 202
68 202
1 6 7 0 0 4224 0 7 6 0 0 2
133 62
116 62
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 240 10
176 79 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 2 0
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
5 4 0.309148 0.500000
344 175 457 272
42991634 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 18 158 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 PWM
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7168 0 0
2
43296 2
0
13 Logic Switch~
5 202 233 0 1 11
0 5
0
0 0 21360 90
2 0V
11 0 25 8
2 V1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
631 0 0
2
43296 1
0
13 Logic Switch~
5 18 103 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 FB
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9466 0 0
2
43296 0
0
14 Logic Display~
6 237 79 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 G1L
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3266 0 0
2
43296 9
0
14 Logic Display~
6 305 78 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 G1L
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7693 0 0
2
43296 8
0
9 Inverter~
13 69 193 0 2 22
0 6 4
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
3723 0 0
2
43296 7
0
5 4013~
219 151 229 0 6 22
0 5 4 7 6 8 2
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U1B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 1 0
1 U
3440 0 0
2
43296 6
0
5 4013~
219 151 139 0 6 22
0 5 6 7 4 9 3
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U1A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 1 0
1 U
6263 0 0
2
43296 5
0
14 Logic Display~
6 237 27 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 G1H
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4900 0 0
2
43296 4
0
14 Logic Display~
6 305 27 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 G2H
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8783 0 0
2
43296 3
0
13
1 0 2 0 0 12432 0 10 0 0 3 5
305 45
305 51
325 51
325 193
237 193
1 0 3 0 0 12304 0 9 0 0 4 4
237 45
237 51
256 51
256 103
6 1 2 0 0 16 0 7 4 0 0 3
175 193
237 193
237 97
6 1 3 0 0 4240 0 8 5 0 0 3
175 103
305 103
305 96
4 0 4 0 0 12432 0 8 0 0 13 4
151 145
151 149
117 149
117 193
1 0 5 0 0 4112 0 2 0 0 8 2
203 220
203 162
4 0 6 0 0 8336 0 7 0 0 12 4
151 235
151 245
43 245
43 193
1 1 5 0 0 12432 0 7 8 0 0 6
151 172
151 162
203 162
203 72
151 72
151 82
1 0 7 0 0 4112 0 1 0 0 11 2
30 158
104 158
1 0 6 0 0 16 0 3 0 0 12 2
30 103
43 103
3 3 7 0 0 8336 0 8 7 0 0 4
127 121
104 121
104 211
127 211
2 1 6 0 0 16 0 8 6 0 0 4
127 103
43 103
43 193
54 193
2 2 4 0 0 16 0 6 7 0 0 6
90 193
117 193
117 191
117 191
117 193
127 193
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

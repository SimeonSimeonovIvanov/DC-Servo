CircuitMaker Text
5.6
Probes: 1
U2_6
Transient Analysis
0 418 47 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 150 10
176 83 1022 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 179 1190 496
9961490 0
0
6 Title:
5 Name:
0
0
0
17
9 Schottky~
219 178 125 0 2 5
0 3 5
0
0 0 848 180
6 11DQ03
-22 -18 20 -10
2 D2
-8 -28 6 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 26108892
68 0 0 0 1 0 0 0
1 D
7978 0 0
2
41826.7 0
0
9 Schottky~
219 248 49 0 2 5
0 4 3
0
0 0 848 180
6 11DQ03
-22 -18 20 -10
2 D1
-8 -28 6 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 26180116
68 0 0 0 1 0 0 0
1 D
3142 0 0
2
41826.7 1
0
10 Op-Amp5:A~
219 172 49 0 5 11
0 2 5 11 12 3
0
0 0 848 0
5 LM358
15 -25 50 -17
2 U1
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 0 0 0
1 U
3284 0 0
2
5.89668e-315 0
0
2 +V
167 172 82 0 1 3
0 12
0
0 0 53616 180
4 -15V
-12 1 16 9
2 V3
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
659 0 0
2
5.89668e-315 5.26354e-315
0
2 +V
167 172 21 0 1 3
0 11
0
0 0 53616 0
4 +15V
-12 -13 16 -5
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3800 0 0
2
5.89668e-315 5.30499e-315
0
7 Ground~
168 145 42 0 1 3
0 2
0
0 0 53360 270
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6792 0 0
2
5.89668e-315 5.32571e-315
0
11 Signal Gen~
195 27 60 0 64 64
0 6 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1092616192
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 1000 0 10 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
7 -10/10V
-25 -30 24 -22
2 V1
-7 -40 7 -32
0
0
37 %D %1 %2 DC 0 SIN(0 10 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3701 0 0
2
5.89668e-315 5.34643e-315
0
7 Ground~
168 69 82 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6316 0 0
2
5.89668e-315 5.3568e-315
0
7 Ground~
168 352 36 0 1 3
0 2
0
0 0 53360 270
0
4 GND3
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8734 0 0
2
5.89668e-315 5.36716e-315
0
2 +V
167 381 15 0 1 3
0 9
0
0 0 53616 0
4 +15V
-12 -13 16 -5
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7988 0 0
2
5.89668e-315 5.37752e-315
0
2 +V
167 381 81 0 1 3
0 10
0
0 0 53616 180
4 -15V
-12 1 16 9
2 V5
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3217 0 0
2
5.89668e-315 5.38788e-315
0
10 Op-Amp5:A~
219 381 43 0 5 11
0 2 7 9 10 8
0
0 0 848 0
5 LM358
15 -25 50 -17
2 U2
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 0 0 0
1 U
3965 0 0
2
5.89668e-315 5.39306e-315
0
11 Resistor:A~
219 115 55 0 2 5
0 6 5
0
0 0 880 0
3 10k
-15 16 6 24
2 R1
-12 6 2 14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8239 0 0
2
5.89668e-315 5.39824e-315
0
11 Resistor:A~
219 213 157 0 2 5
0 5 4
0
0 0 880 0
3 10k
-15 6 6 14
2 R2
-11 -14 3 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
828 0 0
2
5.89668e-315 5.40342e-315
0
11 Resistor:A~
219 385 111 0 2 5
0 7 8
0
0 0 880 0
4 6.8k
-18 6 10 14
2 R5
-11 -14 3 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6187 0 0
2
5.89668e-315 5.4086e-315
0
11 Resistor:A~
219 317 49 0 2 5
0 4 7
0
0 0 880 0
3 10k
-15 16 6 24
2 R3
-12 6 2 14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7107 0 0
2
5.89668e-315 5.41378e-315
0
11 Resistor:A~
219 317 111 0 2 5
0 6 7
0
0 0 880 0
3 20k
-15 6 6 14
2 R4
-11 -14 3 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6433 0 0
2
5.89668e-315 5.41896e-315
0
20
1 1 2 0 0 4096 0 6 3 0 0 2
152 43
154 43
1 0 3 0 0 8320 0 1 0 0 5 3
187 125
219 125
219 49
2 0 4 0 0 8320 0 14 0 0 7 3
231 157
274 157
274 49
2 0 5 0 0 4096 0 1 0 0 17 2
164 125
142 125
2 5 3 0 0 0 0 2 3 0 0 2
234 49
190 49
0 1 6 0 0 8320 0 0 17 16 0 5
82 55
82 185
286 185
286 111
299 111
1 1 4 0 0 0 0 16 2 0 0 2
299 49
257 49
2 0 7 0 0 4096 0 17 0 0 11 2
335 111
349 111
5 2 8 0 0 8320 0 12 15 0 0 4
399 43
419 43
419 111
403 111
1 1 2 0 0 4096 0 9 12 0 0 2
359 37
363 37
1 0 7 0 0 8320 0 15 0 0 14 3
367 111
349 111
349 49
1 3 9 0 0 4224 0 10 12 0 0 2
381 24
381 30
1 4 10 0 0 4224 0 11 12 0 0 2
381 66
381 56
2 2 7 0 0 0 0 16 12 0 0 2
335 49
363 49
1 2 2 0 0 4224 0 8 7 0 0 3
69 76
69 65
58 65
1 1 6 0 0 0 0 7 13 0 0 2
58 55
97 55
1 0 5 0 0 8320 0 14 0 0 20 3
195 157
142 157
142 55
1 3 11 0 0 4224 0 5 3 0 0 2
172 30
172 36
1 4 12 0 0 4224 0 4 3 0 0 2
172 67
172 62
2 2 5 0 0 0 0 13 3 0 0 2
133 55
154 55
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

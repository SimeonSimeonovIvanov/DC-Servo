CircuitMaker Text
5.6
Probes: 1
U3_6
Transient Analysis
0 259 245 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 130 10
176 79 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 2 1
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.563830 0.500000
344 175 2086 704
9961490 0
0
6 Title:
5 Name:
0
0
0
16
10 Op-Amp5:A~
219 230 211 0 5 11
0 9 11 4 3 12
0
0 0 848 0
5 TL082
15 -25 50 -17
2 U3
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 0 0 0
1 U
5433 0 0
2
5.8967e-315 0
0
7 Ground~
168 136 271 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3679 0 0
2
5.8967e-315 0
0
7 Ground~
168 89 144 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9342 0 0
2
43873.9 0
0
11 Signal Gen~
195 33 48 0 64 64
0 7 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1056964608 0 1094713344
0 814313567 814313567 1065353216 1073741824 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 0.5 0 12 0 1e-09 1e-09 1 2 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 0/12V
-18 -30 17 -22
2 FB
-7 -40 7 -32
0
0
37 %D %1 %2 DC 0 PULSE(0 12 0 1n 1n 1 2)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3623 0 0
2
43873.9 1
0
7 Ground~
168 187 101 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3722 0 0
2
43873.9 2
0
14 Opto Isolator~
173 140 55 0 4 9
0 8 10 9 2
0
0 0 880 0
6 OP4N25
-19 19 23 27
2 U1
-22 -27 -8 -19
0
0
17 %D %1 %2 %3 %4 %S
0
0
4 DIP6
9

0 1 2 5 4 1 2 5 4 0
88 0 0 0 1 0 0 0
1 U
8993 0 0
2
43873.9 3
0
14 Opto Isolator~
173 140 120 0 4 9
0 10 2 2 9
0
0 0 880 0
6 OP4N25
-19 19 23 27
2 U2
-22 -27 -8 -19
0
0
17 %D %1 %2 %3 %4 %S
0
0
4 DIP6
9

0 1 2 5 4 1 2 5 4 0
88 0 0 0 1 0 0 0
1 U
3723 0 0
2
43873.9 4
0
11 Signal Gen~
195 33 216 0 64 64
0 6 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1073741824 1084227584 1084227584
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 2 5 5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 0/10V
-18 -30 17 -22
2 SP
-7 -40 7 -32
0
0
35 %D %1 %2 DC 0 SIN(5 5 2 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
6244 0 0
2
43873.9 5
0
7 Ground~
168 100 271 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6421 0 0
2
43873.9 6
0
2 +V
167 230 189 0 1 3
0 4
0
0 0 53616 0
4 +15V
-12 -14 16 -6
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7743 0 0
2
43873.9 7
0
2 +V
167 230 240 0 1 3
0 3
0
0 0 53616 180
4 -15V
-14 0 14 8
2 V5
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9840 0 0
2
43873.9 8
0
11 Resistor:A~
219 136 241 0 3 5
0 2 6 -1
0
0 0 880 90
3 10k
-28 1 -7 9
2 R2
-24 -11 -10 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6910 0 0
2
5.8967e-315 0
0
11 Resistor:A~
219 89 43 0 2 5
0 8 7
0
0 0 880 180
3 560
-11 -14 10 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
449 0 0
2
43873.9 9
0
11 Resistor:A~
219 173 217 0 2 5
0 6 11
0
0 0 880 0
3 51k
-11 18 10 26
2 R4
-7 7 7 15
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8761 0 0
2
43873.9 10
0
11 Resistor:A~
219 173 205 0 2 5
0 6 9
0
0 0 880 0
3 51k
-10 -14 11 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6748 0 0
2
43873.9 11
0
11 Resistor:A~
219 231 271 0 2 5
0 11 12
0
0 0 880 0
3 51k
-12 9 9 17
2 R5
-8 -15 6 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7393 0 0
2
43873.9 12
0
21
4 1 3 0 0 4224 0 1 11 0 0 2
230 224
230 225
3 1 4 0 0 0 0 1 10 0 0 2
230 198
230 198
0 0 5 0 0 0 0 0 0 0 0 2
271 211
271 211
1 1 2 0 0 4096 0 2 12 0 0 2
136 265
136 259
2 0 6 0 0 4096 0 12 0 0 8 2
136 223
136 211
1 0 2 0 0 0 0 3 0 0 7 2
89 138
89 132
2 2 2 0 0 8320 0 7 4 0 0 4
112 132
89 132
89 53
64 53
1 0 6 0 0 4224 0 8 0 0 9 2
64 211
147 211
1 1 6 0 0 0 0 14 15 0 0 4
155 217
147 217
147 205
155 205
1 0 2 0 0 0 0 5 0 0 14 3
187 95
187 87
173 87
1 2 7 0 0 4224 0 4 13 0 0 2
64 43
71 43
1 1 8 0 0 4224 0 13 6 0 0 2
107 43
112 43
0 0 9 0 0 4096 0 0 0 20 15 2
201 205
201 132
4 3 2 0 0 0 0 6 7 0 0 4
166 67
173 67
173 108
166 108
4 3 9 0 0 8320 0 7 6 0 0 4
166 132
201 132
201 43
166 43
1 2 10 0 0 8320 0 7 6 0 0 4
112 108
104 108
104 67
112 67
1 2 2 0 0 0 0 9 8 0 0 3
100 265
100 221
64 221
1 0 11 0 0 8320 0 16 0 0 21 3
213 271
201 271
201 217
5 2 12 0 0 8320 0 1 16 0 0 4
248 211
261 211
261 271
249 271
2 1 9 0 0 0 0 15 1 0 0 2
191 205
212 205
2 2 11 0 0 0 0 14 1 0 0 2
191 217
212 217
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 10 0.002 0.002
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

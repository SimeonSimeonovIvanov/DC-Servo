CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 160 10
176 83 1022 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 2 0
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 179 457 276
42991634 0
0
6 Title:
5 Name:
0
0
0
15
13 Logic Switch~
5 118 226 0 1 11
0 9
0
0 0 21360 90
2 0V
11 0 25 8
2 V1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89666e-315 5.41896e-315
0
13 Logic Switch~
5 26 45 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
7 DIRECTI
-23 -26 26 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89666e-315 5.41378e-315
0
13 Logic Switch~
5 26 100 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 PWM
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89666e-315 5.4086e-315
0
13 Logic Switch~
5 26 154 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
5 BRAKE
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.89666e-315 5.40342e-315
0
14 Logic Display~
6 358 65 0 1 2
10 3
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 G2H
25 0 46 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8157 0 0
2
5.89666e-315 5.39824e-315
0
14 Logic Display~
6 358 8 0 1 2
10 4
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 G1H
25 2 46 10
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
5.89666e-315 5.39306e-315
0
14 Logic Display~
6 358 150 0 1 2
10 5
0
0 0 53872 270
6 100MEG
3 -16 45 -8
6 BREAKE
17 1 59 9
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
5.89666e-315 5.38788e-315
0
5 4013~
219 119 81 0 6 22
0 9 7 8 9 12 13
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U1A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 0 2 1 1 0
1 U
7361 0 0
2
5.89666e-315 5.37752e-315
0
5 4013~
219 119 190 0 6 22
0 9 6 8 9 2 5
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U1B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 0 2 2 1 0
1 U
4747 0 0
2
5.89666e-315 5.36716e-315
0
10 2-In NAND~
219 218 34 0 3 22
0 13 2 4
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
972 0 0
2
5.89666e-315 5.3568e-315
0
10 2-In NAND~
219 218 90 0 3 22
0 12 2 3
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3472 0 0
2
5.89666e-315 5.34643e-315
0
10 2-In NAND~
219 307 43 0 3 22
0 4 2 11
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
9998 0 0
2
5.89666e-315 5.32571e-315
0
10 2-In NAND~
219 306 99 0 3 22
0 3 2 10
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3536 0 0
2
5.89666e-315 5.30499e-315
0
14 Logic Display~
6 358 39 0 1 2
10 11
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 G1L
25 1 46 9
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4597 0 0
2
5.89666e-315 5.26354e-315
0
14 Logic Display~
6 358 95 0 1 2
10 10
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 G2L
25 1 46 9
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3835 0 0
2
5.89666e-315 0
0
21
0 0 2 0 0 4224 0 0 0 17 2 3
180 172
257 172
257 108
2 2 2 0 0 0 0 12 13 0 0 4
283 52
257 52
257 108
282 108
1 0 3 0 0 4224 0 5 0 0 13 3
342 69
273 69
273 90
1 0 4 0 0 4224 0 6 0 0 14 3
342 12
273 12
273 34
1 6 5 0 0 4224 0 7 9 0 0 2
342 154
143 154
1 2 6 0 0 4224 0 4 9 0 0 2
38 154
95 154
1 2 7 0 0 4224 0 2 8 0 0 2
38 45
95 45
1 0 8 0 0 4096 0 3 0 0 9 2
38 100
68 100
3 3 8 0 0 8320 0 9 8 0 0 4
95 172
68 172
68 63
95 63
1 0 9 0 0 4096 0 1 0 0 19 2
119 213
119 204
1 3 10 0 0 4224 0 15 13 0 0 2
342 99
333 99
1 3 11 0 0 4224 0 14 12 0 0 2
342 43
334 43
1 3 3 0 0 0 0 13 11 0 0 2
282 90
245 90
1 3 4 0 0 0 0 12 10 0 0 2
283 34
245 34
1 5 12 0 0 4224 0 11 8 0 0 4
194 81
167 81
167 63
149 63
1 6 13 0 0 4224 0 10 8 0 0 4
194 25
167 25
167 45
143 45
5 0 2 0 0 0 0 9 0 0 18 3
149 172
180 172
180 99
2 2 2 0 0 0 0 10 11 0 0 4
194 43
180 43
180 99
194 99
0 4 9 0 0 4224 0 0 9 21 0 4
83 99
83 204
119 204
119 196
4 0 9 0 0 0 0 8 0 0 21 2
119 87
119 99
1 1 9 0 0 0 0 8 9 0 0 6
119 24
119 11
83 11
83 99
119 99
119 133
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

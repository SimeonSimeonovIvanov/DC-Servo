CircuitMaker Text
5.6
Probes: 1
D2_K
Transient Analysis
0 424 161 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 90 10
176 78 1678 999
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 174 1846 634
9961490 0
0
6 Title:
5 Name:
0
0
0
55
2 +V
167 240 488 0 1 3
0 8
0
0 0 53616 692
4 -15V
-14 1 14 9
2 V8
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3566 0 0
2
41673.5 0
0
7 Ground~
168 265 478 0 1 3
0 2
0
0 0 53360 512
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3371 0 0
2
41673.5 1
0
2 +V
167 240 436 0 1 3
0 9
0
0 0 53616 512
4 +15V
-14 -14 14 -6
3 V13
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4395 0 0
2
41673.5 2
0
8 Op-Amp5~
219 240 460 0 5 11
0 2 6 9 8 7
0
0 0 848 512
5 LM358
-46 -13 -11 -5
3 U3B
-45 -24 -24 -16
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 5 6 8 4 7 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 2 2 0
1 U
6822 0 0
2
41673.5 3
0
2 +V
167 265 346 0 1 3
0 12
0
0 0 53616 90
3 +2V
-10 -16 11 -8
3 V11
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8953 0 0
2
41673.5 4
0
2 +V
167 337 358 0 1 3
0 13
0
0 0 53616 90
5 +2.5V
-42 -5 -7 3
3 V10
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4635 0 0
2
41673.5 5
0
2 +V
167 373 320 0 1 3
0 14
0
0 0 53616 0
4 +15V
-13 -14 15 -6
2 V9
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6596 0 0
2
41673.5 6
0
7 Ground~
168 373 377 0 1 3
0 2
0
0 0 53360 0
0
5 GND15
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3813 0 0
2
41673.5 7
0
8 Op-Amp5~
219 373 350 0 5 11
0 13 11 14 2 10
0
0 0 848 0
5 LM358
15 -25 50 -17
3 U3A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 2 0
1 U
5639 0 0
2
41673.5 8
0
10 Capacitor~
219 573 204 0 2 5
0 5 3
0
0 0 848 692
4 50nF
-11 -19 17 -11
2 C3
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
429 0 0
2
41673.5 9
0
8 Op-Amp5~
219 544 312 0 5 11
0 16 4 17 18 3
0
0 0 848 0
5 LM358
15 -25 50 -17
3 U1B
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 5 6 8 4 7 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 2 1 0
1 U
5832 0 0
2
41673.5 10
0
2 +V
167 544 285 0 1 3
0 17
0
0 0 53616 0
4 +15V
-14 -17 14 -9
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8856 0 0
2
41673.5 11
0
7 Ground~
168 503 377 0 1 3
0 2
0
0 0 53360 0
0
5 GND13
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
469 0 0
2
41673.5 12
0
2 +V
167 544 346 0 1 3
0 18
0
0 0 53616 180
4 -15V
7 -7 35 1
3 V12
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4529 0 0
2
41673.5 13
0
7 Ground~
168 18 333 0 1 3
0 2
0
0 0 53360 512
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
88 0 0
2
5.89649e-315 0
0
7 Ground~
168 83 333 0 1 3
0 2
0
0 0 53360 512
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3894 0 0
2
5.89649e-315 5.26354e-315
0
2 +V
167 83 269 0 1 3
0 25
0
0 0 53616 512
4 +15V
-13 -16 15 -8
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6890 0 0
2
5.89649e-315 5.30499e-315
0
12 Comparator6~
219 85 302 0 6 13
0 7 19 25 2 23 2
0
0 0 848 512
5 LM111
16 -24 51 -16
2 U2
24 -35 38 -27
0
0
23 %D %1 %2 %3 %4 %5 %6 %S
0
0
4 DIP8
13

0 2 3 8 4 7 1 2 3 8
4 7 1 0
88 0 0 256 1 0 0 0
1 U
3257 0 0
2
5.89649e-315 5.32571e-315
0
7 Ground~
168 187 225 0 1 3
0 2
0
0 0 53360 512
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6612 0 0
2
5.89649e-315 5.34643e-315
0
7 Ground~
168 402 225 0 1 3
0 2
0
0 0 53360 512
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3556 0 0
2
5.89649e-315 5.3568e-315
0
7 Ground~
168 117 225 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9143 0 0
2
5.89649e-315 5.36716e-315
0
7 Ground~
168 83 225 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8186 0 0
2
5.89649e-315 5.37752e-315
0
9 Schottky~
219 82 139 0 2 5
0 2 22
0
0 0 848 90
6 1N6392
-53 0 -11 8
2 D1
-52 -12 -38 -4
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
3754 0 0
2
5.89649e-315 5.38788e-315
0
2 +V
167 286 125 0 1 3
0 31
0
0 0 53616 512
4 +15V
-13 -15 15 -7
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8708 0 0
2
5.89649e-315 5.39306e-315
0
7 Ground~
168 373 225 0 1 3
0 2
0
0 0 53360 512
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3338 0 0
2
5.89649e-315 5.39824e-315
0
8 Op-Amp5~
219 286 161 0 5 11
0 28 29 31 2 30
0
0 0 848 0
5 LM358
7 -16 42 -8
3 U1A
8 -25 29 -17
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 1 0
1 U
5546 0 0
2
5.89649e-315 5.40342e-315
0
7 Ground~
168 250 225 0 1 3
0 2
0
0 0 53360 512
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3295 0 0
2
5.89649e-315 5.4086e-315
0
12 Zener Diode~
219 373 194 0 2 5
0 2 15
0
0 0 848 602
6 1N4731
-59 -1 -17 7
2 D2
-57 -13 -43 -5
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
100 0 0 0 1 0 0 0
1 D
4923 0 0
2
5.89649e-315 5.41378e-315
0
7 Ground~
168 286 225 0 1 3
0 2
0
0 0 53360 512
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3248 0 0
2
5.89649e-315 5.41896e-315
0
10 Capacitor~
219 187 195 0 2 5
0 27 2
0
0 0 848 782
4 10nF
13 6 41 14
2 C2
12 -4 26 4
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3139 0 0
2
5.89649e-315 5.42414e-315
0
9 Inductor~
219 117 139 0 2 5
0 22 26
0
0 0 848 270
3 2mH
12 -1 33 7
2 L1
12 -11 26 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
3285 0 0
2
5.89649e-315 5.42933e-315
0
2 +V
167 19 20 0 1 3
0 21
0
0 0 53616 512
4 +25V
-13 -14 15 -6
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
336 0 0
2
5.89649e-315 5.43192e-315
0
12 PNP Trans:C~
219 78 83 0 3 7
0 22 24 21
0
0 0 848 692
7 FZT792A
17 0 66 8
2 Q1
35 -10 49 -2
0
0
14 %D %1 %2 %3 %M
0
0
7 SOT-223
7

0 2 1 3 2 1 3 0
113 0 0 0 1 0 0 0
1 Q
6582 0 0
2
5.89649e-315 5.43451e-315
0
2 +V
167 82 373 0 1 3
0 20
0
0 0 53616 512
3 +5V
-11 -13 10 -5
2 V7
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3546 0 0
2
5.89649e-315 5.4371e-315
0
7 Ground~
168 82 478 0 1 3
0 2
0
0 0 53360 512
0
5 GND12
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
893 0 0
2
5.89649e-315 5.43969e-315
0
7 Ground~
168 118 478 0 1 3
0 2
0
0 0 53360 512
0
5 GND11
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8998 0 0
2
5.89649e-315 5.44228e-315
0
4 VCO~
221 109 425 0 5 9
0 20 2 19 2 3
0
0 0 80 0
6 TRIVCO
37 -2 79 6
2 V6
36 -2 50 6
0
0
29 %D %%vd(%1,%2) %%vd(%3,%4) %M
0
96 alias:ATRIVCO {LOW=0 HIGH=5 CYCLE=0.000255 C1=5 C2=0 C3=0 C4=0 C5=0 F1=4000 F2=0 F3=0 F4=0 F5=0}
0
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 V
5979 0 0
2
5.89649e-315 5.44487e-315
0
11 Resistor:A~
219 221 411 0 2 5
0 6 7
0
0 0 880 512
2 1k
-14 -16 0 -8
3 R13
-13 -26 8 -18
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3835 0 0
2
41673.5 14
0
11 Resistor:A~
219 310 411 0 2 5
0 6 3
0
0 0 880 692
2 1k
-16 -15 -2 -7
3 R15
-15 -24 6 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
750 0 0
2
41673.5 15
0
11 Resistor:A~
219 368 292 0 2 5
0 11 10
0
0 0 880 0
2 1k
-7 -14 7 -6
3 R18
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
849 0 0
2
41673.5 16
0
11 Resistor:A~
219 306 344 0 4 5
0 11 12 0 1
0
0 0 880 180
2 1k
-7 -14 7 -6
3 R16
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4693 0 0
2
41673.5 17
0
11 Resistor:A~
219 534 204 0 2 5
0 4 5
0
0 0 880 0
2 1K
-8 -14 6 -6
3 R14
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4775 0 0
2
41673.5 18
0
11 Resistor:A~
219 468 205 0 2 5
0 4 10
0
0 0 880 180
3 10k
-11 -14 10 -6
3 R17
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9572 0 0
2
41673.5 19
0
11 Resistor:A~
219 546 161 0 2 5
0 4 3
0
0 0 880 0
4 9.5k
-13 -14 15 -6
3 R12
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3761 0 0
2
41673.5 20
0
11 Resistor:A~
219 467 161 0 2 5
0 4 15
0
0 0 880 180
3 10k
-11 -14 10 -6
3 R11
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6765 0 0
2
41673.5 21
0
11 Resistor:A~
219 503 345 0 3 5
0 2 16 -1
0
0 0 880 90
2 1k
11 0 25 8
3 R10
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7938 0 0
2
41673.5 22
0
11 Resistor:A~
219 19 192 0 2 5
0 24 23
0
0 0 880 782
4 2.7k
9 -1 37 7
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
55 0 0
2
5.89649e-315 5.44746e-315
0
11 Resistor:A~
219 216 167 0 2 5
0 28 27
0
0 0 880 512
2 1k
-12 8 2 16
2 R5
-13 -14 1 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5610 0 0
2
5.89649e-315 5.45005e-315
0
11 Resistor:A~
219 158 167 0 2 5
0 27 26
0
0 0 880 512
2 1k
-12 7 2 15
2 R4
-12 -15 2 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3322 0 0
2
5.89649e-315 5.45264e-315
0
9 Resistor~
219 117 193 0 3 5
0 2 26 -1
0
0 0 880 90
3 0.1
5 0 26 8
2 R3
6 -11 20 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5914 0 0
2
5.89649e-315 5.45523e-315
0
11 Resistor:A~
219 250 196 0 3 5
0 2 29 -1
0
0 0 880 602
2 2k
8 2 22 10
2 R6
8 -9 22 -1
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8748 0 0
2
5.89649e-315 5.45782e-315
0
11 Resistor:A~
219 343 103 0 2 5
0 29 15
0
0 0 880 692
3 18K
-10 -14 11 -6
2 R7
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5830 0 0
2
5.89649e-315 5.46041e-315
0
11 Resistor:A~
219 343 161 0 2 5
0 30 15
0
0 0 880 692
2 1K
-7 -14 7 -6
2 R8
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9153 0 0
2
5.89649e-315 5.463e-315
0
9 Resistor~
219 402 193 0 3 5
0 2 15 -1
0
0 0 880 602
2 1k
8 0 22 8
2 R9
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9220 0 0
2
5.89649e-315 5.46559e-315
0
11 Resistor:A~
219 19 57 0 3 5
0 21 24 1
0
0 0 880 782
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7901 0 0
2
5.89649e-315 5.46818e-315
0
61
2 0 3 0 0 4224 0 39 0 0 5 3
328 411
604 411
604 312
2 0 3 0 0 0 0 44 0 0 5 3
564 161
604 161
604 204
0 0 4 0 0 4096 0 0 0 6 4 2
503 205
503 161
1 1 4 0 0 0 0 45 44 0 0 2
485 161
528 161
2 5 3 0 0 0 0 10 11 0 0 4
582 204
604 204
604 312
562 312
2 0 4 0 0 8320 0 11 0 0 8 3
526 306
503 306
503 205
1 2 5 0 0 4224 0 10 42 0 0 2
564 204
552 204
1 1 4 0 0 0 0 42 43 0 0 3
516 204
516 205
486 205
1 0 6 0 0 4096 0 39 0 0 10 2
292 411
265 411
1 2 6 0 0 8320 0 38 4 0 0 4
239 411
265 411
265 454
258 454
1 0 7 0 0 8320 0 18 0 0 14 3
101 308
179 308
179 411
1 4 8 0 0 0 0 1 4 0 0 2
240 473
240 473
1 1 2 0 0 8192 0 2 4 0 0 3
265 472
265 466
258 466
5 2 7 0 0 0 0 4 38 0 0 4
222 460
179 460
179 411
203 411
1 3 9 0 0 4224 0 3 4 0 0 2
240 445
240 447
2 0 10 0 0 8320 0 43 0 0 17 3
450 205
427 205
427 292
2 5 10 0 0 0 0 40 9 0 0 4
386 292
427 292
427 350
391 350
1 0 11 0 0 8320 0 40 0 0 20 3
350 292
338 292
338 344
1 2 12 0 0 4224 0 5 41 0 0 2
276 344
288 344
1 2 11 0 0 0 0 41 9 0 0 2
324 344
355 344
1 1 13 0 0 4224 0 6 9 0 0 2
348 356
355 356
1 3 14 0 0 4224 0 7 9 0 0 2
373 329
373 337
1 4 2 0 0 4096 0 8 9 0 0 2
373 371
373 363
2 0 15 0 0 4096 0 45 0 0 54 2
449 161
402 161
2 1 16 0 0 8320 0 46 11 0 0 3
503 327
503 318
526 318
1 1 2 0 0 0 0 46 13 0 0 2
503 363
503 371
1 3 17 0 0 4224 0 12 11 0 0 2
544 294
544 299
1 4 18 0 0 4224 0 14 11 0 0 2
544 331
544 325
3 2 19 0 0 4224 0 37 18 0 0 3
118 401
118 296
101 296
1 4 2 0 0 4096 0 36 37 0 0 2
118 472
118 455
1 2 2 0 0 0 0 35 37 0 0 2
82 472
82 455
1 1 20 0 0 4224 0 37 34 0 0 2
82 401
82 382
0 3 21 0 0 4224 0 0 33 40 0 3
19 35
83 35
83 65
1 6 2 0 0 8192 0 15 18 0 0 3
18 327
18 310
67 310
1 4 2 0 0 0 0 16 18 0 0 2
83 327
83 315
1 0 22 0 0 8320 0 31 0 0 43 3
117 121
117 112
83 112
2 5 23 0 0 4224 0 47 18 0 0 3
19 210
19 294
67 294
2 0 24 0 0 4096 0 33 0 0 39 2
60 83
19 83
2 1 24 0 0 4224 0 55 47 0 0 2
19 75
19 174
1 1 21 0 0 0 0 32 55 0 0 2
19 29
19 39
1 3 25 0 0 4224 0 17 18 0 0 2
83 278
83 289
2 0 26 0 0 4224 0 49 0 0 46 2
140 167
117 167
2 1 22 0 0 0 0 23 33 0 0 2
83 126
83 101
1 1 2 0 0 4224 0 22 23 0 0 2
83 219
83 149
1 1 2 0 0 0 0 21 50 0 0 2
117 219
117 211
2 2 26 0 0 0 0 50 31 0 0 2
117 175
117 157
2 1 2 0 0 0 0 30 19 0 0 2
187 204
187 219
1 0 27 0 0 4096 0 30 0 0 49 2
187 186
187 167
1 2 27 0 0 4224 0 49 48 0 0 2
176 167
198 167
1 1 28 0 0 4224 0 48 26 0 0 2
234 167
268 167
2 0 29 0 0 4096 0 51 0 0 53 2
250 178
250 155
2 0 15 0 0 8320 0 52 0 0 54 3
361 103
373 103
373 161
1 2 29 0 0 4224 0 52 26 0 0 4
325 103
250 103
250 155
268 155
2 0 15 0 0 0 0 54 0 0 58 3
402 175
402 161
373 161
1 1 2 0 0 0 0 20 54 0 0 2
402 219
402 211
1 4 2 0 0 0 0 29 26 0 0 2
286 219
286 174
1 1 2 0 0 0 0 25 28 0 0 2
373 219
373 204
2 2 15 0 0 0 0 28 53 0 0 3
373 184
373 161
361 161
1 5 30 0 0 4224 0 53 26 0 0 4
325 161
303 161
303 161
304 161
1 1 2 0 0 0 0 27 51 0 0 2
250 219
250 214
1 3 31 0 0 4224 0 24 26 0 0 2
286 134
286 148
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
226 289 308 313
230 294 303 310
11 SP Current:
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.02 1e-06 1e-06
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

CircuitMaker Text
5.6
Probes: 1
U1B_7
Transient Analysis
0 509 171 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 130 10
176 79 1918 540
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 2 0
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
2 2 0.500000 0.500000
344 175 2086 645
9961490 0
0
6 Title:
5 Name:
0
0
0
45
12 Zener Diode~
219 391 10 0 2 5
0 32 4
0
0 0 848 180
7 1N4745A
-26 -22 23 -14
2 D4
-9 -32 5 -24
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 26094748
100 0 0 768 1 1 0 0
1 D
7699 0 0
2
43873.9 0
0
12 Zener Diode~
219 438 10 0 2 5
0 33 5
0
0 0 848 0
7 1N4745A
-22 -22 27 -14
2 D3
-5 -32 9 -24
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 26211368
100 0 0 768 1 1 0 0
1 D
6638 0 0
2
43873.9 1
0
10 Capacitor~
219 415 63 0 2 5
0 4 3
0
0 0 848 0
5 3.3nF
-17 -18 18 -10
2 C3
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4595 0 0
2
43873.9 2
0
7 Ground~
168 1038 319 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9395 0 0
2
5.89668e-315 0
0
10 Capacitor~
219 446 102 0 2 5
0 20 5
0
0 0 848 0
5 100nF
-19 -18 16 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3303 0 0
2
5.89668e-315 5.26354e-315
0
8 Op-Amp5~
219 412 173 0 5 11
0 2 4 23 22 3
0
0 0 848 0
5 TL082
15 -25 50 -17
3 U1B
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 5 6 8 4 7 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 2 1 0
1 U
4498 0 0
2
5.89668e-315 5.30499e-315
0
8 Op-Amp5~
219 217 167 0 5 11
0 2 29 25 24 28
0
0 0 848 0
5 TL082
15 -25 50 -17
3 U1A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 1 0
1 U
9728 0 0
2
5.89668e-315 5.32571e-315
0
7 Ground~
168 117 298 0 1 3
0 2
0
0 0 53360 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3789 0 0
2
5.89668e-315 5.34643e-315
0
11 Signal Gen~
195 52 264 0 64 64
0 27 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1101004800 -1054867456 1092616192
0 814313567 814313567 1020054733 1028443341 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 20 -10 10 0 1e-09 1e-09 0.025 0.05 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
7 -10/10V
-25 -30 24 -22
2 V7
-7 -40 7 -32
0
0
43 %D %1 %2 DC 0 PULSE(-10 10 0 1n 1n 25m 50m)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3978 0 0
2
5.89668e-315 5.3568e-315
0
7 Ground~
168 444 284 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3494 0 0
2
5.89668e-315 5.36716e-315
0
14 Var ResistorA~
219 448 205 0 3 7
0 21 5 3
0
0 0 848 602
7 10k 10%
3 4 52 12
3 R11
6 -13 27 -5
0
0
30 %DA %1 %2 1000
%DB %2 %3 9000
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
82 0 0 0 1 0 0 0
1 R
3507 0 0
2
5.89668e-315 5.37752e-315
0
7 Ground~
168 379 285 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5151 0 0
2
5.89668e-315 5.38788e-315
0
2 +V
167 412 150 0 1 3
0 23
0
0 0 53616 0
4 +15V
-14 -13 14 -5
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3701 0 0
2
5.89668e-315 5.39306e-315
0
2 +V
167 412 201 0 1 3
0 22
0
0 0 53616 180
4 -15V
-13 -1 15 7
2 V3
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8585 0 0
2
5.89668e-315 5.39824e-315
0
2 +V
167 217 195 0 1 3
0 24
0
0 0 53616 180
4 -15V
-13 -1 15 7
2 V2
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8809 0 0
2
5.89668e-315 5.40342e-315
0
2 +V
167 217 144 0 1 3
0 25
0
0 0 53616 0
4 +15V
-14 -13 14 -5
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5993 0 0
2
5.89668e-315 5.4086e-315
0
7 Ground~
168 189 190 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8654 0 0
2
5.89668e-315 5.41378e-315
0
7 Ground~
168 60 190 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7223 0 0
2
5.89668e-315 5.41896e-315
0
14 Var ResistorA~
219 64 163 0 3 7
0 2 30 31
0
0 0 848 602
7 10k 80%
-61 -4 -12 4
2 R2
-43 -14 -29 -6
0
0
30 %DA %1 %2 8000
%DB %2 %3 2000
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
82 0 0 0 1 0 0 0
1 R
3641 0 0
2
5.89668e-315 5.42414e-315
0
8 Op-Amp5~
219 786 173 0 5 11
0 2 8 16 15 11
0
0 0 848 0
5 TL082
15 -25 50 -17
3 U2A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 2 0
1 U
3104 0 0
2
5.89668e-315 5.42933e-315
0
10 Capacitor~
219 949 126 0 2 5
0 12 7
0
0 0 848 0
6 1000nF
-23 -19 19 -11
2 C2
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3296 0 0
2
5.89668e-315 5.43192e-315
0
2 +V
167 786 206 0 1 3
0 15
0
0 0 53616 180
5 -100V
-16 -1 19 7
2 V8
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8534 0 0
2
5.89668e-315 5.43451e-315
0
2 +V
167 786 147 0 1 3
0 16
0
0 0 53616 0
5 +100V
-17 -13 18 -5
2 V9
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
949 0 0
2
5.89668e-315 5.4371e-315
0
7 Ground~
168 756 196 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3371 0 0
2
5.89668e-315 5.43969e-315
0
7 Ground~
168 869 203 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7311 0 0
2
5.89668e-315 5.44228e-315
0
2 +V
167 946 158 0 1 3
0 14
0
0 0 53616 0
4 100V
-14 -13 14 -5
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3409 0 0
2
5.89668e-315 5.44487e-315
0
2 +V
167 946 210 0 1 3
0 13
0
0 0 53616 180
5 -100V
-17 -2 18 6
2 V6
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3526 0 0
2
5.89668e-315 5.44746e-315
0
8 Op-Amp5~
219 946 181 0 5 11
0 11 12 14 13 7
0
0 0 848 0
5 TL082
15 -25 50 -17
3 U2B
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 5 6 8 4 7 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 2 2 0
1 U
4129 0 0
2
5.89668e-315 5.45005e-315
0
8 Op-Amp5~
219 645 167 0 5 11
0 10 9 19 18 9
0
0 0 848 0
5 TL082
15 -25 50 -17
3 U3A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 3 0
1 U
6278 0 0
2
5.89668e-315 5.45264e-315
0
2 +V
167 645 144 0 1 3
0 19
0
0 0 53616 0
4 +15V
-14 -13 14 -5
3 V11
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3482 0 0
2
5.89668e-315 5.45523e-315
0
2 +V
167 645 195 0 1 3
0 18
0
0 0 53616 180
4 -15V
-13 -1 15 7
3 V10
7 -12 28 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8323 0 0
2
5.89668e-315 5.45782e-315
0
11 Resistor:A~
219 1038 281 0 3 5
0 2 6 -1
0
0 0 880 90
2 1k
10 0 24 8
3 R18
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3984 0 0
2
5.89668e-315 5.46041e-315
0
11 Resistor:A~
219 1038 215 0 2 5
0 6 7
0
0 0 880 90
2 9k
10 0 24 8
3 R17
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7622 0 0
2
5.89668e-315 5.463e-315
0
11 Resistor:A~
219 393 102 0 2 5
0 4 20
0
0 0 880 0
4 500k
-14 -14 14 -6
3 R10
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
816 0 0
2
5.89668e-315 5.46559e-315
0
11 Resistor:A~
219 444 246 0 3 5
0 2 21 -1
0
0 0 880 90
3 15k
6 0 27 8
2 R6
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4656 0 0
2
5.89668e-315 5.46818e-315
0
11 Resistor:A~
219 320 167 0 2 5
0 28 4
0
0 0 880 0
3 20k
-10 -14 11 -6
2 R8
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6356 0 0
2
5.89668e-315 5.47077e-315
0
11 Resistor:A~
219 157 102 0 2 5
0 27 29
0
0 0 880 0
4 220k
-13 -14 15 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7479 0 0
2
5.89668e-315 5.47207e-315
0
11 Resistor:A~
219 222 102 0 2 5
0 29 28
0
0 0 880 0
4 220k
-13 -14 15 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5690 0 0
2
5.89668e-315 5.47336e-315
0
11 Resistor:A~
219 157 161 0 2 5
0 30 29
0
0 0 880 0
4 220k
-13 -14 15 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5617 0 0
2
5.89668e-315 5.47466e-315
0
11 Resistor:A~
219 60 105 0 2 5
0 31 7
0
0 0 880 90
3 15k
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3903 0 0
2
5.89668e-315 5.47595e-315
0
11 Resistor:A~
219 800 123 0 2 5
0 8 11
0
0 0 880 0
4 100k
-13 -14 15 -6
3 R13
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4452 0 0
2
5.89668e-315 5.47725e-315
0
11 Resistor:A~
219 728 167 0 2 5
0 9 8
0
0 0 880 0
3 10k
-10 -14 11 -6
3 R14
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6282 0 0
2
5.89668e-315 5.47854e-315
0
11 Resistor:A~
219 900 175 0 3 5
0 2 12 -1
0
0 0 880 0
3 10k
-10 -14 11 -6
3 R12
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7187 0 0
2
5.89668e-315 5.47984e-315
0
11 Resistor:A~
219 538 173 0 2 5
0 3 17
0
0 0 880 0
3 10k
-10 -14 11 -6
3 R16
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6866 0 0
2
5.89668e-315 5.48113e-315
0
11 Resistor:A~
219 588 173 0 2 5
0 17 10
0
0 0 880 0
3 10k
-10 -14 11 -6
3 R15
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7670 0 0
2
5.89668e-315 5.48243e-315
0
53
2 0 3 0 0 8320 0 3 0 0 14 3
424 63
501 63
501 173
1 0 4 0 0 4096 0 3 0 0 5 2
406 63
352 63
0 1 4 0 0 0 0 0 3 0 0 2
406 63
406 63
2 0 5 0 0 8192 0 2 0 0 31 3
448 10
482 10
482 102
0 2 4 0 0 4224 0 0 1 32 0 3
352 102
352 10
381 10
1 1 2 0 0 4096 0 10 35 0 0 2
444 278
444 264
1 1 2 0 0 0 0 4 32 0 0 2
1038 313
1038 299
2 1 6 0 0 4224 0 32 33 0 0 2
1038 263
1038 233
2 0 7 0 0 4096 0 33 0 0 30 2
1038 197
1038 181
1 0 8 0 0 8320 0 41 0 0 11 3
782 123
756 123
756 167
2 2 8 0 0 0 0 20 42 0 0 2
768 167
746 167
1 0 9 0 0 4096 0 42 0 0 27 2
710 167
699 167
1 2 10 0 0 4224 0 29 45 0 0 2
627 173
606 173
1 0 3 0 0 0 0 44 0 0 42 2
520 173
444 173
2 0 11 0 0 8192 0 41 0 0 16 3
818 123
839 123
839 187
1 5 11 0 0 4224 0 28 20 0 0 4
928 187
824 187
824 173
804 173
2 5 7 0 0 4096 0 21 28 0 0 4
958 126
1014 126
1014 181
964 181
1 0 12 0 0 8320 0 21 0 0 22 3
940 126
922 126
922 175
1 1 2 0 0 4096 0 25 43 0 0 3
869 197
869 175
882 175
4 1 13 0 0 4224 0 28 27 0 0 2
946 194
946 195
3 1 14 0 0 4224 0 28 26 0 0 2
946 168
946 167
2 2 12 0 0 0 0 43 28 0 0 2
918 175
928 175
4 1 15 0 0 4224 0 20 22 0 0 2
786 186
786 191
3 1 16 0 0 4224 0 20 23 0 0 2
786 160
786 156
1 1 2 0 0 0 0 24 20 0 0 3
756 190
756 179
768 179
2 1 17 0 0 4224 0 44 45 0 0 2
556 173
570 173
2 5 9 0 0 12416 0 29 29 0 0 6
627 161
617 161
617 125
699 125
699 167
663 167
4 1 18 0 0 0 0 29 31 0 0 2
645 180
645 180
3 1 19 0 0 4224 0 29 30 0 0 2
645 154
645 153
2 0 7 0 0 8320 0 40 0 0 17 5
60 87
60 29
1038 29
1038 181
1014 181
2 2 5 0 0 8320 0 11 5 0 0 4
456 203
482 203
482 102
455 102
1 0 4 0 0 0 0 34 0 0 45 3
375 102
352 102
352 167
2 1 20 0 0 4224 0 34 5 0 0 2
411 102
437 102
2 1 21 0 0 4224 0 35 11 0 0 2
444 228
444 219
4 1 22 0 0 0 0 6 14 0 0 2
412 186
412 186
3 1 23 0 0 4224 0 6 13 0 0 2
412 160
412 159
4 1 24 0 0 0 0 7 15 0 0 2
217 180
217 180
3 1 25 0 0 4224 0 7 16 0 0 2
217 154
217 153
0 0 26 0 0 0 0 0 0 0 0 2
854 4
854 4
1 2 2 0 0 8192 0 8 9 0 0 3
117 292
117 269
83 269
1 1 27 0 0 8320 0 9 37 0 0 4
83 259
116 259
116 102
139 102
3 5 3 0 0 0 0 11 6 0 0 3
444 183
444 173
430 173
1 2 28 0 0 4096 0 36 0 0 51 2
302 167
266 167
1 1 2 0 0 4224 0 12 6 0 0 3
379 279
379 179
394 179
2 2 4 0 0 0 0 6 36 0 0 2
394 167
338 167
2 0 29 0 0 4096 0 37 0 0 47 2
175 102
189 102
1 0 29 0 0 8320 0 38 0 0 50 3
204 102
189 102
189 161
1 2 30 0 0 4224 0 39 19 0 0 2
139 161
72 161
1 1 2 0 0 0 0 17 7 0 0 3
189 184
189 173
199 173
2 2 29 0 0 0 0 7 39 0 0 2
199 161
175 161
2 5 28 0 0 8320 0 38 7 0 0 4
240 102
266 102
266 167
235 167
1 1 2 0 0 0 0 18 19 0 0 2
60 184
60 177
3 1 31 0 0 4224 0 19 40 0 0 2
60 141
60 123
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.25 0.0001 0.0001
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

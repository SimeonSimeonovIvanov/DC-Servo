CircuitMaker Text
5.6
Probes: 1
C1_2
Transient Analysis
0 467 97 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 160 10
176 79 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 2 0
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 457 272
9961490 0
0
6 Title:
5 Name:
0
0
0
25
8 Op-Amp5~
219 189 91 0 5 11
0 14 15 17 16 12
0
0 0 832 0
5 TL082
8 -15 43 -7
3 U1A
15 -26 36 -18
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 1 0
1 U
5130 0 0
2
43283 0
0
2 +V
167 189 68 0 1 3
0 17
0
0 0 53600 0
4 +15V
-14 -14 14 -6
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
391 0 0
2
43283 1
0
2 +V
167 189 120 0 1 3
0 16
0
0 0 53600 180
4 -15V
-12 -1 16 7
2 V2
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3124 0 0
2
43283 2
0
7 Ground~
168 117 162 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3421 0 0
2
43283 3
0
7 Ground~
168 154 162 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8157 0 0
2
43283 4
0
11 Signal Gen~
195 29 90 0 64 64
0 13 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1036831949 -1054867456 1092616192
0 814313567 814313567 1084227584 1092616192 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 26
20
0 0.1 -10 10 0 1e-09 1e-09 5 10 0
0 0 0 0 0 0 0 0 0 0
0
0 0 1344 0
7 -10/10V
-25 -30 24 -22
2 V5
-7 -40 7 -32
8 Speed SP
-27 -40 29 -32
0
40 %D %1 %2 DC 0 PULSE(-10 10 0 1n 1n 5 10)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
5572 0 0
2
43283 5
0
7 Ground~
168 87 162 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8901 0 0
2
43283 6
0
6 Diode~
219 261 91 0 2 5
0 12 10
0
0 0 832 0
6 1N4148
-21 -18 21 -10
2 D2
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
7361 0 0
2
43283 7
0
6 Diode~
219 261 44 0 2 5
0 11 12
0
0 0 832 180
6 1N4148
-21 -18 21 -10
2 D1
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
4747 0 0
2
43283 8
0
14 Var ResistorA~
219 310 52 0 3 7
0 3 3 11
0
0 0 832 180
7 5k7 50%
-22 -25 27 -17
3 RP1
-9 -36 12 -28
0
0
30 %DA %1 %2 2500
%DB %2 %3 2500
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
82 0 0 0 1 0 0 0
1 R
972 0 0
2
43283 9
0
14 Var ResistorA~
219 310 91 0 3 7
0 3 3 10
0
0 0 832 512
8 5k7 0.1%
-29 18 27 26
3 RP2
-10 8 11 16
0
0
27 %DA %1 %2 5
%DB %2 %3 4995
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
82 0 0 0 1 0 0 0
1 R
3472 0 0
2
43283 10
0
7 Ground~
168 343 162 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9998 0 0
2
43283 11
0
10 Capacitor~
219 465 44 0 2 5
0 7 5
0
0 0 832 0
3 1uF
-12 -18 9 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3536 0 0
2
43283 12
0
2 +V
167 428 74 0 1 3
0 8
0
0 0 53600 0
4 +15V
-14 -14 14 -6
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4597 0 0
2
43283 13
0
2 +V
167 428 126 0 1 3
0 9
0
0 0 53600 180
4 -15V
-12 -1 16 7
2 V3
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3835 0 0
2
43283 14
0
7 Ground~
168 402 162 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3670 0 0
2
43283 15
0
8 Op-Amp5~
219 428 97 0 5 11
0 4 6 8 9 5
0
0 0 832 0
5 TL082
10 -14 45 -6
3 U1B
16 -25 37 -17
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 5 6 8 4 7 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 2 1 0
1 U
5616 0 0
2
43283 16
0
11 Resistor:A~
219 402 129 0 4 5
0 4 2 0 -1
0
0 0 864 270
3 10k
-29 1 -8 9
2 R8
-25 -11 -11 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9323 0 0
2
43283 17
0
11 Resistor:A~
219 427 44 0 2 5
0 7 6
0
0 0 864 180
5 0.001
-16 -14 19 -6
2 R7
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
317 0 0
2
43283 18
0
11 Resistor:A~
219 89 85 0 2 5
0 15 13
0
0 0 864 180
4 1.3k
-14 -14 14 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3108 0 0
2
43283 19
0
11 Resistor:A~
219 117 128 0 3 5
0 2 15 -1
0
0 0 864 90
3 10k
-27 0 -6 8
2 R2
-24 -10 -10 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4299 0 0
2
43283 20
0
11 Resistor:A~
219 154 54 0 2 5
0 14 5
0
0 0 864 90
4 1.3k
-35 1 -7 9
2 R3
-29 -8 -15 0
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9672 0 0
2
43283 21
0
11 Resistor:A~
219 154 128 0 3 5
0 2 14 -1
0
0 0 864 90
3 10k
-28 -1 -7 7
2 R4
-24 -11 -10 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7876 0 0
2
43283 22
0
11 Resistor:A~
219 343 128 0 4 5
0 3 2 0 -1
0
0 0 864 270
4 1.3k
-39 4 -11 12
2 R5
-31 -6 -17 2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6369 0 0
2
43283 23
0
11 Resistor:A~
219 372 91 0 2 5
0 6 3
0
0 0 864 180
4 220k
-13 -14 15 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9172 0 0
2
43283 24
0
29
2 0 3 0 0 4096 0 25 0 0 13 2
354 91
343 91
1 1 4 0 0 4224 0 18 17 0 0 3
402 111
402 103
410 103
2 1 2 0 0 4096 0 18 16 0 0 2
402 147
402 156
2 0 3 0 0 8192 0 11 0 0 14 3
312 79
312 71
343 71
2 0 3 0 0 0 0 10 0 0 14 3
312 56
312 64
343 64
0 2 5 0 0 8320 0 0 22 10 0 4
484 44
484 4
154 4
154 36
2 0 6 0 0 8320 0 19 0 0 9 3
409 44
402 44
402 91
1 1 7 0 0 4224 0 19 13 0 0 2
445 44
456 44
1 2 6 0 0 0 0 25 17 0 0 2
390 91
410 91
2 5 5 0 0 0 0 13 17 0 0 4
474 44
484 44
484 97
446 97
1 3 8 0 0 4224 0 14 17 0 0 2
428 83
428 84
1 4 9 0 0 4224 0 15 17 0 0 2
428 111
428 110
1 0 3 0 0 0 0 24 0 0 14 2
343 110
343 91
1 1 3 0 0 8320 0 10 11 0 0 4
328 44
343 44
343 91
328 91
3 2 10 0 0 4224 0 11 8 0 0 2
292 91
271 91
3 1 11 0 0 4224 0 10 9 0 0 2
292 44
271 44
1 0 12 0 0 4096 0 8 0 0 18 2
251 91
237 91
2 5 12 0 0 8320 0 9 1 0 0 4
251 44
237 44
237 91
207 91
1 2 2 0 0 4096 0 12 24 0 0 2
343 156
343 146
2 1 2 0 0 8320 0 6 7 0 0 3
60 95
87 95
87 156
1 2 13 0 0 4224 0 6 20 0 0 2
60 85
71 85
1 1 2 0 0 0 0 5 23 0 0 2
154 156
154 146
1 1 2 0 0 0 0 4 21 0 0 2
117 156
117 146
1 0 14 0 0 4096 0 1 0 0 25 2
171 97
154 97
2 1 14 0 0 4224 0 23 22 0 0 2
154 110
154 72
2 0 15 0 0 4096 0 21 0 0 27 2
117 110
117 85
1 2 15 0 0 4224 0 20 1 0 0 2
107 85
171 85
1 4 16 0 0 4224 0 3 1 0 0 2
189 105
189 104
1 3 17 0 0 4224 0 2 1 0 0 2
189 77
189 78
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 50 0.02 0.02
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

CircuitMaker Text
5.6
Probes: 1
D2_K
Transient Analysis
0 363 119 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 210 10
176 83 1022 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 2 1
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 179 1190 496
9961490 0
0
6 Title:
5 Name:
0
0
0
19
7 Ground~
168 95 165 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8239 0 0
2
5.89682e-315 5.41896e-315
0
8 Op-Amp5~
219 122 92 0 5 11
0 15 14 17 16 8
0
0 0 848 0
5 TL082
15 -25 50 -17
3 U1A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 0 2 1 1 0
1 U
828 0 0
2
5.89682e-315 5.41378e-315
0
2 +V
167 122 120 0 1 3
0 16
0
0 0 53616 180
4 -15V
-14 0 14 8
2 V1
-7 -10 7 -2
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6187 0 0
2
5.89682e-315 5.4086e-315
0
2 +V
167 122 70 0 1 3
0 17
0
0 0 53616 0
4 +15V
-13 -14 15 -6
2 V2
-6 -24 8 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7107 0 0
2
5.89682e-315 5.40342e-315
0
2 +V
167 198 94 0 1 3
0 7
0
0 0 54640 90
5 -0.5V
-16 5 19 13
2 V3
-6 -5 8 3
5 TACHO
-15 -17 20 -9
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6433 0 0
2
5.89682e-315 5.39824e-315
0
2 +V
167 11 88 0 1 3
0 9
0
0 0 54640 90
2 2V
-4 5 10 13
2 V4
-4 -3 10 5
2 SP
-4 -16 10 -8
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8559 0 0
2
5.89682e-315 5.39306e-315
0
2 +V
167 253 30 0 1 3
0 13
0
0 0 53616 0
4 +15V
-13 -14 15 -6
2 V5
-6 -24 8 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3674 0 0
2
5.89682e-315 5.38788e-315
0
2 +V
167 253 80 0 1 3
0 12
0
0 0 53616 180
4 -15V
-14 0 14 8
2 V6
-7 -10 7 -2
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5697 0 0
2
5.89682e-315 5.37752e-315
0
8 Op-Amp5~
219 253 52 0 5 11
0 7 9 13 12 5
0
0 0 848 0
5 TL082
15 -25 50 -17
3 U1B
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 5 6 8 4 7 3 2 8 4
1 5 6 8 4 7 0
88 0 0 0 2 2 1 0
1 U
3805 0 0
2
5.89682e-315 5.36716e-315
0
8 Op-Amp5~
219 253 135 0 5 11
0 8 7 11 10 6
0
0 0 848 0
5 TL082
15 -25 50 -17
3 U2A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 0 2 1 2 0
1 U
5219 0 0
2
5.89682e-315 5.3568e-315
0
2 +V
167 253 163 0 1 3
0 10
0
0 0 53616 180
4 -15V
-14 0 14 8
2 V7
-7 -10 7 -2
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3795 0 0
2
5.89682e-315 5.34643e-315
0
2 +V
167 253 113 0 1 3
0 11
0
0 0 53616 0
4 +15V
-13 -14 15 -6
2 V8
-6 -24 8 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3637 0 0
2
5.89682e-315 5.32571e-315
0
6 Diode~
219 329 52 0 2 5
0 5 4
0
0 0 848 0
6 1N4148
-21 -18 21 -10
2 D1
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
3226 0 0
2
5.89682e-315 5.30499e-315
0
6 Diode~
219 331 135 0 2 5
0 6 4
0
0 0 848 0
6 1N4148
-21 -18 21 -10
2 D2
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
6966 0 0
2
5.89682e-315 5.26354e-315
0
2 +V
167 363 209 0 1 3
0 3
0
0 0 53616 180
4 -15V
-14 0 14 8
2 V9
-7 -10 7 -2
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9796 0 0
2
5.89682e-315 0
0
11 Resistor:A~
219 95 133 0 4 5
0 15 2 0 -1
0
0 0 880 270
4 5.1k
-35 -2 -7 6
2 R1
-28 -12 -14 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5952 0 0
2
5.89682e-315 5.43451e-315
0
11 Resistor:A~
219 123 46 0 2 5
0 8 14
0
0 0 880 180
3 10k
-11 -14 10 -6
2 R2
-8 -24 6 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3649 0 0
2
5.89682e-315 5.43192e-315
0
11 Resistor:A~
219 67 86 0 4 5
0 14 9 0 1
0
0 0 880 180
3 10k
-11 -14 10 -6
2 R3
-8 -24 6 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3716 0 0
2
5.89682e-315 5.42933e-315
0
11 Resistor:A~
219 363 166 0 4 5
0 4 3 0 1
0
0 0 880 270
3 15k
-32 -2 -11 6
2 R4
-29 -12 -15 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4797 0 0
2
5.89682e-315 5.42414e-315
0
21
1 2 3 0 0 4224 0 15 19 0 0 2
363 194
363 184
1 0 4 0 0 4096 0 19 0 0 3 2
363 148
363 135
2 2 4 0 0 8320 0 13 14 0 0 4
339 52
363 52
363 135
341 135
5 1 5 0 0 4224 0 9 13 0 0 2
271 52
319 52
1 5 6 0 0 4224 0 14 10 0 0 2
321 135
271 135
1 0 7 0 0 4096 0 5 0 0 7 2
209 92
225 92
2 1 7 0 0 8320 0 10 9 0 0 4
235 129
225 129
225 58
235 58
1 0 8 0 0 4224 0 10 0 0 15 3
235 141
173 141
173 91
2 0 9 0 0 12416 0 9 0 0 14 5
235 46
225 46
225 1
38 1
38 86
1 4 10 0 0 0 0 11 10 0 0 2
253 148
253 148
1 3 11 0 0 0 0 12 10 0 0 2
253 122
253 122
1 4 12 0 0 0 0 8 9 0 0 2
253 65
253 65
1 3 13 0 0 0 0 7 9 0 0 2
253 39
253 39
1 2 9 0 0 0 0 6 18 0 0 2
22 86
49 86
1 5 8 0 0 0 0 17 2 0 0 4
141 46
173 46
173 92
140 92
2 1 2 0 0 4224 0 16 1 0 0 2
95 151
95 159
2 0 14 0 0 8320 0 17 0 0 21 3
105 46
95 46
95 86
1 1 15 0 0 4224 0 16 2 0 0 3
95 115
95 98
104 98
1 4 16 0 0 0 0 3 2 0 0 2
122 105
122 105
1 3 17 0 0 0 0 4 2 0 0 2
122 79
122 79
1 2 14 0 0 0 0 18 2 0 0 2
85 86
104 86
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

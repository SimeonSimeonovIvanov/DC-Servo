CircuitMaker Text
5.6
Probes: 1
D2_K
Transient Analysis
0 405 163 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 150 10
176 78 1678 999
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.272530 0.500000
344 174 1846 425
9961490 0
0
6 Title:
5 Name:
0
0
0
85
8 Op-Amp5~
219 871 329 0 5 11
0 9 8 10 11 4
0
0 0 848 0
5 LM358
15 -25 50 -17
3 U6A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 5 0
1 U
4382 0 0
2
41673.5 3
0
2 +V
167 871 302 0 1 3
0 10
0
0 0 53616 0
4 +15V
-14 -17 14 -9
3 V12
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4748 0 0
2
41673.5 2
0
7 Ground~
168 830 394 0 1 3
0 2
0
0 0 53360 0
0
5 GND13
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7459 0 0
2
41673.5 1
0
2 +V
167 871 363 0 1 3
0 11
0
0 0 53616 180
4 -15V
7 -7 35 1
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9955 0 0
2
41673.5 0
0
8 Op-Amp5~
219 696 483 0 5 11
0 15 14 16 17 5
0
0 0 848 0
5 LM358
12 -11 47 -3
3 U5B
12 -23 33 -15
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 5 6 8 4 7 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 2 4 0
1 U
3116 0 0
2
41673.5 25
0
2 +V
167 696 456 0 1 3
0 16
0
0 0 53616 0
4 +15V
-15 -14 13 -6
3 V20
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7963 0 0
2
41673.5 24
0
7 Ground~
168 661 548 0 1 3
0 2
0
0 0 53360 0
0
5 GND18
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9310 0 0
2
41673.5 23
0
2 +V
167 696 517 0 1 3
0 17
0
0 0 53616 180
4 -15V
-12 0 16 8
3 V19
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8679 0 0
2
41673.5 22
0
8 Op-Amp5~
219 696 167 0 5 11
0 19 18 20 21 6
0
0 0 848 0
5 LM358
14 -11 49 -3
3 U5A
14 -23 35 -15
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 4 0
1 U
6856 0 0
2
41673.5 21
0
2 +V
167 696 140 0 1 3
0 20
0
0 0 53616 0
4 +15V
-14 -14 14 -6
3 V18
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
333 0 0
2
41673.5 20
0
7 Ground~
168 661 232 0 1 3
0 2
0
0 0 53360 0
0
5 GND17
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7356 0 0
2
41673.5 19
0
2 +V
167 696 201 0 1 3
0 21
0
0 0 53616 180
4 -15V
-13 0 15 8
3 V17
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8964 0 0
2
41673.5 18
0
2 +V
167 696 363 0 1 3
0 26
0
0 0 53616 180
4 -15V
-13 -1 15 7
3 V16
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8173 0 0
2
41673.5 17
0
7 Ground~
168 661 394 0 1 3
0 2
0
0 0 53360 0
0
5 GND16
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3349 0 0
2
41673.5 16
0
2 +V
167 696 302 0 1 3
0 25
0
0 0 53616 0
4 +15V
-14 -14 14 -6
3 V15
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9520 0 0
2
41673.5 15
0
8 Op-Amp5~
219 696 329 0 5 11
0 24 22 25 26 7
0
0 0 848 0
5 LM358
14 -11 49 -3
3 U4B
14 -24 35 -16
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 5 6 8 4 7 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 2 3 0
1 U
3112 0 0
2
41673.5 14
0
10 Capacitor~
219 727 272 0 2 5
0 23 7
0
0 0 848 692
4 10nF
-11 -19 17 -11
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3731 0 0
2
41673.5 13
0
10 Capacitor~
219 619 477 0 2 5
0 14 13
0
0 0 848 512
3 1nF
-11 -18 10 -10
2 C3
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6631 0 0
2
41673.5 8
0
2 +V
167 536 248 0 1 3
0 30
0
0 0 53616 180
4 -15V
7 -7 35 1
3 V14
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3802 0 0
2
41673.5 7
0
7 Ground~
168 495 279 0 1 3
0 2
0
0 0 53360 0
0
5 GND14
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5487 0 0
2
41673.5 6
0
2 +V
167 536 187 0 1 3
0 29
0
0 0 53616 0
4 +15V
-14 -17 14 -9
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
672 0 0
2
41673.5 5
0
8 Op-Amp5~
219 536 214 0 5 11
0 28 27 29 30 13
0
0 0 848 0
5 LM358
15 -25 50 -17
3 U4A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 3 0
1 U
5836 0 0
2
41673.5 4
0
7 Ground~
168 400 548 0 1 3
0 2
0
0 0 53360 512
0
5 GND20
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9906 0 0
2
41673.5 0
0
2 +V
167 373 454 0 1 3
0 34
0
0 0 53616 512
4 +15V
-14 -14 14 -6
3 V21
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
891 0 0
2
41673.5 4
0
7 Ground~
168 373 548 0 1 3
0 2
0
0 0 53360 512
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3694 0 0
2
41673.5 3
0
8 Op-Amp5~
219 373 483 0 5 11
0 33 32 34 2 31
0
0 0 848 512
5 LM358
-45 -15 -10 -7
3 U6B
-44 -27 -23 -19
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 5 6 8 4 7 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 2 5 0
1 U
5372 0 0
2
41673.5 2
0
2 +V
167 265 346 0 1 3
0 36
0
0 0 53616 90
3 +2V
-10 -16 11 -8
3 V11
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5178 0 0
2
41673.5 4
0
2 +V
167 337 358 0 1 3
0 37
0
0 0 53616 90
5 +2.5V
-42 -5 -7 3
3 V10
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
514 0 0
2
41673.5 5
0
2 +V
167 373 320 0 1 3
0 38
0
0 0 53616 0
4 +15V
-13 -14 15 -6
2 V9
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3447 0 0
2
41673.5 6
0
7 Ground~
168 373 377 0 1 3
0 2
0
0 0 53360 0
0
5 GND15
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4800 0 0
2
41673.5 7
0
8 Op-Amp5~
219 373 350 0 5 11
0 37 35 38 2 12
0
0 0 848 0
5 LM358
15 -25 50 -17
3 U3A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 2 0
1 U
9835 0 0
2
41673.5 8
0
7 Ground~
168 18 333 0 1 3
0 2
0
0 0 53360 512
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5194 0 0
2
5.89649e-315 0
0
7 Ground~
168 83 333 0 1 3
0 2
0
0 0 53360 512
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3807 0 0
2
5.89649e-315 5.26354e-315
0
2 +V
167 83 269 0 1 3
0 45
0
0 0 53616 512
4 +15V
-13 -16 15 -8
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3650 0 0
2
5.89649e-315 5.30499e-315
0
12 Comparator6~
219 85 302 0 6 13
0 31 39 45 2 43 2
0
0 0 848 512
5 LM111
16 -24 51 -16
2 U2
24 -35 38 -27
0
0
23 %D %1 %2 %3 %4 %5 %6 %S
0
0
4 DIP8
13

0 2 3 8 4 7 1 2 3 8
4 7 1 0
88 0 0 256 1 0 0 0
1 U
4310 0 0
2
5.89649e-315 5.32571e-315
0
7 Ground~
168 187 225 0 1 3
0 2
0
0 0 53360 512
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4278 0 0
2
5.89649e-315 5.34643e-315
0
7 Ground~
168 402 225 0 1 3
0 2
0
0 0 53360 512
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
765 0 0
2
5.89649e-315 5.3568e-315
0
7 Ground~
168 117 225 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7128 0 0
2
5.89649e-315 5.36716e-315
0
7 Ground~
168 83 225 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
374 0 0
2
5.89649e-315 5.37752e-315
0
9 Schottky~
219 82 139 0 2 5
0 2 42
0
0 0 848 90
6 1N6392
-53 0 -11 8
2 D1
-52 -12 -38 -4
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
6381 0 0
2
5.89649e-315 5.38788e-315
0
2 +V
167 286 125 0 1 3
0 51
0
0 0 53616 512
4 +15V
-13 -15 15 -7
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3410 0 0
2
5.89649e-315 5.39306e-315
0
7 Ground~
168 373 225 0 1 3
0 2
0
0 0 53360 512
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7522 0 0
2
5.89649e-315 5.39824e-315
0
8 Op-Amp5~
219 286 161 0 5 11
0 48 49 51 2 50
0
0 0 848 0
5 LM358
7 -16 42 -8
3 U1A
8 -25 29 -17
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 1 0
1 U
8978 0 0
2
5.89649e-315 5.40342e-315
0
7 Ground~
168 250 225 0 1 3
0 2
0
0 0 53360 512
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7148 0 0
2
5.89649e-315 5.4086e-315
0
12 Zener Diode~
219 373 194 0 2 5
0 2 3
0
0 0 848 602
6 1N4731
-59 -1 -17 7
2 D2
-57 -13 -43 -5
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
100 0 0 0 1 0 0 0
1 D
9514 0 0
2
5.89649e-315 5.41378e-315
0
7 Ground~
168 286 225 0 1 3
0 2
0
0 0 53360 512
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3720 0 0
2
5.89649e-315 5.41896e-315
0
10 Capacitor~
219 187 195 0 2 5
0 47 2
0
0 0 848 782
4 10nF
13 6 41 14
2 C2
12 -4 26 4
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
489 0 0
2
5.89649e-315 5.42414e-315
0
9 Inductor~
219 117 139 0 2 5
0 42 46
0
0 0 848 270
3 1mH
12 -1 33 7
2 L1
12 -11 26 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
3307 0 0
2
5.89649e-315 5.42933e-315
0
2 +V
167 19 20 0 1 3
0 41
0
0 0 53616 512
4 +50V
-13 -14 15 -6
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8816 0 0
2
5.89649e-315 5.43192e-315
0
12 PNP Trans:C~
219 78 83 0 3 7
0 42 44 41
0
0 0 848 692
7 FZT792A
17 0 66 8
2 Q1
35 -10 49 -2
0
0
14 %D %1 %2 %3 %M
0
0
7 SOT-223
7

0 2 1 3 2 1 3 0
113 0 0 0 1 0 0 0
1 Q
3809 0 0
2
5.89649e-315 5.43451e-315
0
2 +V
167 82 373 0 1 3
0 40
0
0 0 53616 512
3 +5V
-11 -13 10 -5
2 V7
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5816 0 0
2
5.89649e-315 5.4371e-315
0
7 Ground~
168 82 478 0 1 3
0 2
0
0 0 53360 512
0
5 GND12
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8733 0 0
2
5.89649e-315 5.43969e-315
0
7 Ground~
168 118 478 0 1 3
0 2
0
0 0 53360 512
0
5 GND11
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5111 0 0
2
5.89649e-315 5.44228e-315
0
4 VCO~
221 109 425 0 5 9
0 40 2 39 2 3
0
0 0 80 0
6 TRIVCO
37 -2 79 6
2 V6
36 -2 50 6
0
0
29 %D %%vd(%1,%2) %%vd(%3,%4) %M
0
96 alias:ATRIVCO {LOW=0 HIGH=5 CYCLE=0.000255 C1=5 C2=0 C3=0 C4=0 C5=0 F1=4000 F2=0 F3=0 F4=0 F5=0}
0
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 V
3992 0 0
2
5.89649e-315 5.44487e-315
0
11 Resistor:A~
219 799 323 0 2 5
0 8 5
0
0 0 880 180
3 10k
-11 -14 10 -6
3 R32
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5751 0 0
2
41673.5 8
0
11 Resistor:A~
219 799 261 0 2 5
0 8 6
0
0 0 880 180
3 10k
-11 -14 10 -6
3 R17
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9211 0 0
2
41673.5 7
0
11 Resistor:A~
219 873 261 0 2 5
0 8 4
0
0 0 880 0
3 10k
-10 -14 11 -6
3 R14
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8222 0 0
2
41673.5 6
0
11 Resistor:A~
219 799 292 0 2 5
0 8 7
0
0 0 880 180
6 10000k
-21 -14 21 -6
3 R12
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3198 0 0
2
41673.5 5
0
11 Resistor:A~
219 830 362 0 3 5
0 2 9 -1
0
0 0 880 90
2 1k
-29 1 -15 9
3 R11
-30 -11 -9 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4605 0 0
2
41673.5 4
0
11 Resistor:A~
219 661 516 0 3 5
0 2 15 -1
0
0 0 880 90
2 1k
-29 1 -15 9
3 R29
-30 -11 -9 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8683 0 0
2
41673.5 38
0
11 Resistor:A~
219 703 114 0 2 5
0 18 6
0
0 0 880 0
3 10k
-10 -14 11 -6
3 R28
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3998 0 0
2
41673.5 37
0
11 Resistor:A~
219 620 161 0 2 5
0 18 13
0
0 0 880 180
3 10k
-11 -14 10 -6
3 R27
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3778 0 0
2
41673.5 36
0
11 Resistor:A~
219 661 200 0 3 5
0 2 19 -1
0
0 0 880 90
2 1k
-29 1 -15 9
3 R26
-30 -11 -9 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7433 0 0
2
41673.5 35
0
11 Resistor:A~
219 619 323 0 2 5
0 22 13
0
0 0 880 180
2 5k
-8 -14 6 -6
3 R24
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3224 0 0
2
41673.5 34
0
11 Resistor:A~
219 661 362 0 3 5
0 2 24 -1
0
0 0 880 90
2 1k
-26 0 -12 8
3 R25
-30 -12 -9 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6792 0 0
2
41673.5 33
0
11 Resistor:A~
219 686 272 0 2 5
0 22 23
0
0 0 880 0
1 1
-5 -14 2 -6
3 R19
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5935 0 0
2
41673.5 32
0
11 Resistor:A~
219 704 430 0 2 5
0 14 5
0
0 0 880 0
2 1K
-8 -14 6 -6
3 R30
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6381 0 0
2
41673.5 26
0
11 Resistor:A~
219 495 247 0 3 5
0 2 28 -1
0
0 0 880 90
2 1k
-29 1 -15 9
3 R23
-30 -11 -9 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4685 0 0
2
41673.5 3
0
11 Resistor:A~
219 465 208 0 2 5
0 27 12
0
0 0 880 180
3 10k
-11 -14 10 -6
3 R22
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
346 0 0
2
41673.5 2
0
11 Resistor:A~
219 538 161 0 2 5
0 27 13
0
0 0 880 0
3 10k
-10 -14 11 -6
3 R21
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5219 0 0
2
41673.5 1
0
11 Resistor:A~
219 464 161 0 2 5
0 27 3
0
0 0 880 180
3 10k
-11 -14 10 -6
3 R20
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3107 0 0
2
41673.5 0
0
11 Resistor:A~
219 400 513 0 4 5
0 33 2 0 -1
0
0 0 880 782
2 1k
11 0 25 8
3 R15
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3665 0 0
2
41673.5 0
0
11 Resistor:A~
219 361 427 0 2 5
0 32 31
0
0 0 880 512
2 1k
-7 -14 7 -6
3 R10
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9374 0 0
2
41673.5 1
0
11 Resistor:A~
219 449 477 0 2 5
0 32 4
0
0 0 880 692
2 1k
-7 -14 7 -6
3 R13
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4937 0 0
2
41673.5 0
0
11 Resistor:A~
219 368 292 0 2 5
0 35 12
0
0 0 880 0
2 1k
-7 -14 7 -6
3 R18
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8929 0 0
2
41673.5 16
0
11 Resistor:A~
219 306 344 0 4 5
0 35 36 0 1
0
0 0 880 180
2 1k
-7 -14 7 -6
3 R16
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5165 0 0
2
41673.5 17
0
11 Resistor:A~
219 19 192 0 2 5
0 44 43
0
0 0 880 782
4 2.7k
9 -1 37 7
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9550 0 0
2
5.89649e-315 5.44746e-315
0
11 Resistor:A~
219 216 167 0 2 5
0 48 47
0
0 0 880 512
2 1k
-12 8 2 16
2 R5
-13 -14 1 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6272 0 0
2
5.89649e-315 5.45005e-315
0
11 Resistor:A~
219 158 167 0 2 5
0 47 46
0
0 0 880 512
2 1k
-12 7 2 15
2 R4
-12 -15 2 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7647 0 0
2
5.89649e-315 5.45264e-315
0
9 Resistor~
219 117 193 0 3 5
0 2 46 -1
0
0 0 880 90
3 0.1
5 0 26 8
2 R3
6 -11 20 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4145 0 0
2
5.89649e-315 5.45523e-315
0
11 Resistor:A~
219 250 196 0 3 5
0 2 49 -1
0
0 0 880 602
2 2k
8 2 22 10
2 R6
8 -9 22 -1
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3589 0 0
2
5.89649e-315 5.45782e-315
0
11 Resistor:A~
219 343 103 0 2 5
0 49 3
0
0 0 880 692
3 18K
-10 -14 11 -6
2 R7
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4480 0 0
2
5.89649e-315 5.46041e-315
0
11 Resistor:A~
219 343 161 0 2 5
0 50 3
0
0 0 880 692
2 1K
-7 -14 7 -6
2 R8
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4488 0 0
2
5.89649e-315 5.463e-315
0
9 Resistor~
219 402 193 0 3 5
0 2 3 -1
0
0 0 880 602
3 10k
4 0 25 8
2 R9
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5788 0 0
2
5.89649e-315 5.46559e-315
0
11 Resistor:A~
219 19 57 0 3 5
0 41 44 1
0
0 0 880 782
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3334 0 0
2
5.89649e-315 5.46818e-315
0
96
2 0 3 0 0 4096 0 84 0 0 4 2
402 175
402 161
2 0 3 0 0 4096 0 45 0 0 3 2
373 184
373 161
2 0 3 0 0 8192 0 82 0 0 4 3
361 103
373 103
373 161
2 2 3 0 0 4224 0 71 83 0 0 2
446 161
361 161
2 0 4 0 0 12416 0 74 0 0 12 5
467 477
495 477
495 567
921 567
921 329
2 0 5 0 0 8320 0 55 0 0 23 4
781 323
767 323
767 483
750 483
2 0 6 0 0 8320 0 56 0 0 30 4
781 261
767 261
767 167
751 167
2 0 7 0 0 4096 0 58 0 0 36 2
781 292
752 292
1 0 8 0 0 4096 0 58 0 0 10 2
817 292
830 292
0 0 8 0 0 4224 0 0 0 11 13 2
830 323
830 261
1 2 8 0 0 0 0 55 1 0 0 2
817 323
853 323
5 2 4 0 0 0 0 1 57 0 0 4
889 329
921 329
921 261
891 261
1 1 8 0 0 0 0 56 57 0 0 2
817 261
855 261
2 1 9 0 0 8320 0 59 1 0 0 3
830 344
830 335
853 335
1 1 2 0 0 4096 0 59 3 0 0 2
830 380
830 388
1 3 10 0 0 4224 0 2 1 0 0 2
871 311
871 316
1 4 11 0 0 4224 0 4 1 0 0 2
871 348
871 342
2 0 12 0 0 8320 0 69 0 0 60 3
447 208
427 208
427 292
2 0 13 0 0 4096 0 64 0 0 20 2
601 323
586 323
0 2 13 0 0 4224 0 0 18 44 0 3
586 214
586 477
610 477
2 0 13 0 0 0 0 62 0 0 44 2
602 161
586 161
1 0 14 0 0 8192 0 67 0 0 24 3
686 430
661 430
661 477
5 2 5 0 0 0 0 5 67 0 0 4
714 483
752 483
752 430
722 430
2 1 14 0 0 4224 0 5 18 0 0 2
678 477
628 477
2 1 15 0 0 8320 0 60 5 0 0 3
661 498
661 489
678 489
1 1 2 0 0 0 0 60 7 0 0 2
661 534
661 542
1 3 16 0 0 4224 0 6 5 0 0 2
696 465
696 470
1 4 17 0 0 4224 0 8 5 0 0 2
696 502
696 496
1 0 18 0 0 8320 0 61 0 0 31 3
685 114
661 114
661 161
5 2 6 0 0 0 0 9 61 0 0 4
714 167
752 167
752 114
721 114
2 1 18 0 0 0 0 9 62 0 0 2
678 161
638 161
2 1 19 0 0 8320 0 63 9 0 0 3
661 182
661 173
678 173
1 1 2 0 0 0 0 63 11 0 0 2
661 218
661 226
1 3 20 0 0 4224 0 10 9 0 0 2
696 149
696 154
1 4 21 0 0 4224 0 12 9 0 0 2
696 186
696 180
5 2 7 0 0 8320 0 16 17 0 0 4
714 329
752 329
752 272
736 272
1 0 22 0 0 8320 0 66 0 0 38 3
668 272
661 272
661 323
1 2 22 0 0 0 0 64 16 0 0 2
637 323
678 323
1 2 23 0 0 4224 0 17 66 0 0 2
718 272
704 272
2 1 24 0 0 8320 0 65 16 0 0 3
661 344
661 335
678 335
1 1 2 0 0 0 0 65 14 0 0 2
661 380
661 388
1 3 25 0 0 4224 0 15 16 0 0 2
696 311
696 316
1 4 26 0 0 4224 0 13 16 0 0 2
696 348
696 342
5 2 13 0 0 0 0 22 70 0 0 4
554 214
586 214
586 161
556 161
0 0 27 0 0 4224 0 0 0 47 46 2
495 208
495 161
1 1 27 0 0 0 0 71 70 0 0 2
482 161
520 161
2 1 27 0 0 0 0 22 69 0 0 2
518 208
483 208
2 1 28 0 0 8320 0 68 22 0 0 3
495 229
495 220
518 220
1 1 2 0 0 0 0 68 20 0 0 2
495 265
495 273
1 3 29 0 0 4224 0 21 22 0 0 2
536 196
536 201
1 4 30 0 0 4224 0 19 22 0 0 2
536 233
536 227
0 1 31 0 0 8336 0 0 35 53 0 4
319 483
187 483
187 308
101 308
2 5 31 0 0 0 0 73 26 0 0 4
343 427
319 427
319 483
355 483
1 0 32 0 0 8320 0 73 0 0 59 3
379 427
400 427
400 477
1 2 2 0 0 4096 0 23 72 0 0 2
400 542
400 531
1 1 33 0 0 8320 0 72 26 0 0 3
400 495
400 489
391 489
1 4 2 0 0 4096 0 25 26 0 0 2
373 542
373 496
1 3 34 0 0 4224 0 24 26 0 0 2
373 463
373 470
1 2 32 0 0 0 0 74 26 0 0 6
431 477
400 477
400 476
400 476
400 477
391 477
2 5 12 0 0 0 0 75 31 0 0 4
386 292
427 292
427 350
391 350
1 0 35 0 0 8320 0 75 0 0 63 3
350 292
338 292
338 344
1 2 36 0 0 4224 0 27 76 0 0 2
276 344
288 344
1 2 35 0 0 0 0 76 31 0 0 2
324 344
355 344
1 1 37 0 0 4224 0 28 31 0 0 2
348 356
355 356
1 3 38 0 0 4224 0 29 31 0 0 2
373 329
373 337
1 4 2 0 0 0 0 30 31 0 0 2
373 371
373 363
3 2 39 0 0 4224 0 54 35 0 0 3
118 401
118 296
101 296
1 4 2 0 0 0 0 53 54 0 0 2
118 472
118 455
1 2 2 0 0 0 0 52 54 0 0 2
82 472
82 455
1 1 40 0 0 4224 0 54 51 0 0 2
82 401
82 382
0 3 41 0 0 4224 0 0 50 78 0 3
19 35
83 35
83 65
1 6 2 0 0 8192 0 32 35 0 0 3
18 327
18 310
67 310
1 4 2 0 0 0 0 33 35 0 0 2
83 327
83 315
1 0 42 0 0 8320 0 48 0 0 81 3
117 121
117 112
83 112
2 5 43 0 0 4224 0 77 35 0 0 3
19 210
19 294
67 294
2 0 44 0 0 4096 0 50 0 0 77 2
60 83
19 83
2 1 44 0 0 4224 0 85 77 0 0 2
19 75
19 174
1 1 41 0 0 0 0 49 85 0 0 2
19 29
19 39
1 3 45 0 0 4224 0 34 35 0 0 2
83 278
83 289
2 0 46 0 0 4224 0 79 0 0 84 2
140 167
117 167
2 1 42 0 0 0 0 40 50 0 0 2
83 126
83 101
1 1 2 0 0 4224 0 39 40 0 0 2
83 219
83 149
1 1 2 0 0 0 0 38 80 0 0 2
117 219
117 211
2 2 46 0 0 0 0 80 48 0 0 2
117 175
117 157
2 1 2 0 0 0 0 47 36 0 0 2
187 204
187 219
1 0 47 0 0 4096 0 47 0 0 87 2
187 186
187 167
1 2 47 0 0 4224 0 79 78 0 0 2
176 167
198 167
1 1 48 0 0 4224 0 78 43 0 0 2
234 167
268 167
2 0 49 0 0 4096 0 81 0 0 90 2
250 178
250 155
1 2 49 0 0 4224 0 82 43 0 0 4
325 103
250 103
250 155
268 155
1 1 2 0 0 0 0 37 84 0 0 2
402 219
402 211
1 4 2 0 0 0 0 46 43 0 0 2
286 219
286 174
1 1 2 0 0 0 0 42 45 0 0 2
373 219
373 204
1 5 50 0 0 4224 0 83 43 0 0 4
325 161
303 161
303 161
304 161
1 1 2 0 0 0 0 44 81 0 0 2
250 219
250 214
1 3 51 0 0 4224 0 41 43 0 0 2
286 134
286 148
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
226 289 308 313
230 294 303 310
11 SP Current:
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.02 1e-06 1e-06
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

CircuitMaker Text
5.6
Probes: 1
R1_2
Transient Analysis
0 169 118 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 170 10
427 83 1678 999
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 2 0
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.356987 0.500000
595 179 1846 506
9961490 0
0
6 Title:
5 Name:
0
0
0
24
10 P-EMOS 3T~
219 554 160 0 3 7
0 3 9 11
0
0 0 848 512
7 IRF7104
-71 0 -22 8
2 Q4
-53 -10 -39 -2
0
0
17 %D %1 %2 %3 %3 %M
0
0
16 SMD8A(A:8,1,2)(B
7

0 1 2 3 1 2 3 0
109 0 0 256 0 0 0 0
1 Q
7502 0 0
2
41950.5 23
0
2 +V
167 611 187 0 1 3
0 9
0
0 0 53616 602
4 -15V
-13 -15 15 -7
2 V3
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
7826 0 0
2
41950.5 22
0
7 Ground~
168 544 247 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5360 0 0
2
41950.5 21
0
10 P-EMOS 3T~
219 554 209 0 3 7
0 2 9 11
0
0 0 848 180
7 IRF7104
-71 0 -22 8
2 Q3
-53 -10 -39 -2
0
0
17 %D %1 %2 %3 %3 %M
0
0
16 SMD8A(A:8,1,2)(B
7

0 1 2 3 1 2 3 0
109 0 0 256 0 0 0 0
1 Q
3543 0 0
2
41950.5 20
0
7 Ground~
168 404 248 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4527 0 0
2
41950.5 19
0
14 Var ResistorA~
219 459 53 0 3 7
0 5 12 10
0
0 0 848 90
7 10k 50%
16 -2 65 6
3 R10
24 -16 45 -8
0
0
30 %DA %1 %2 5000
%DB %2 %3 5000
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
82 0 0 0 0 0 0 0
1 R
4230 0 0
2
41950.5 18
0
7 Ground~
168 463 247 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4851 0 0
2
41950.5 17
0
11 Signal Gen~
195 49 191 0 64 64
0 10 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1120403456 0 1050253722
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 22
20
1 100 0 0.3 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
11 -300m/300mV
-39 -30 38 -22
2 V1
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 SIN(0 300m 100 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
3665 0 0
2
41950.5 8
0
7 Ground~
168 94 246 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9874 0 0
2
41950.5 7
0
7 Ground~
168 188 248 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
793 0 0
2
41950.5 6
0
14 Var ResistorA~
219 184 122 0 3 7
0 15 14 8
0
0 0 848 90
7 10k 99%
16 -2 65 6
2 R1
27 -16 41 -8
0
0
29 %DA %1 %2 9900
%DB %2 %3 100
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
82 0 0 0 0 0 0 0
1 R
9424 0 0
2
41950.5 5
0
7 Ground~
168 129 249 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9751 0 0
2
41950.5 4
0
10 P-EMOS 3T~
219 279 210 0 3 7
0 2 9 13
0
0 0 848 180
7 IRF7104
-71 0 -22 8
2 Q1
-53 -10 -39 -2
0
0
17 %D %1 %2 %3 %3 %M
0
0
16 SMD8A(A:8,1,2)(B
7

0 1 2 3 1 2 3 0
109 0 0 256 0 0 0 0
1 Q
6169 0 0
2
41950.5 3
0
7 Ground~
168 269 248 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3362 0 0
2
41950.5 2
0
10 P-EMOS 3T~
219 279 161 0 3 7
0 7 9 13
0
0 0 848 512
7 IRF7104
-71 0 -22 8
2 Q2
-53 -10 -39 -2
0
0
17 %D %1 %2 %3 %3 %M
0
0
16 SMD8A(A:8,1,2)(B
7

0 1 2 3 1 2 3 0
109 0 0 256 0 0 0 0
1 Q
4391 0 0
2
41950.5 0
0
9 Resistor~
219 511 88 0 2 5
0 4 5
0
0 0 880 180
4 2.7k
-14 -14 14 -6
3 R11
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
8214 0 0
2
41950.6 1
0
9 Resistor~
219 544 117 0 2 5
0 3 4
0
0 0 880 90
2 1k
10 0 24 8
2 R8
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
7266 0 0
2
41950.6 0
0
9 Resistor~
219 269 116 0 2 5
0 7 6
0
0 0 880 90
3 10k
6 0 27 8
2 R9
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3947 0 0
2
41950.6 0
0
11 Resistor:A~
219 404 188 0 3 5
0 2 12 -1
0
0 0 880 90
6 10000k
9 2 51 10
2 R7
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
5715 0 0
2
41950.5 14
0
9 Resistor~
219 463 185 0 3 5
0 2 5 -1
0
0 0 880 90
4 5.1k
2 0 30 8
2 R6
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
5703 0 0
2
41950.5 13
0
9 Resistor~
219 188 186 0 3 5
0 2 15 -1
0
0 0 880 90
4 2.7k
2 0 30 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3511 0 0
2
41950.5 12
0
11 Resistor:A~
219 129 189 0 3 5
0 2 14 -1
0
0 0 880 90
6 10000k
9 2 51 10
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9901 0 0
2
41950.5 11
0
9 Resistor~
219 235 88 0 2 5
0 6 8
0
0 0 880 180
4 2.7k
-14 -14 14 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9115 0 0
2
41950.5 10
0
9 Resistor~
219 188 51 0 2 5
0 8 10
0
0 0 880 90
4 5.1k
7 0 35 8
2 R5
13 -10 27 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
5545 0 0
2
41950.5 9
0
26
1 1 3 0 0 4224 0 17 1 0 0 2
544 135
544 142
2 1 4 0 0 8336 0 17 16 0 0 3
544 99
544 88
529 88
2 0 5 0 0 4112 0 16 0 0 15 2
493 88
463 88
2 1 6 0 0 8320 0 18 23 0 0 3
269 98
269 88
253 88
1 1 7 0 0 4224 0 18 15 0 0 2
269 134
269 143
2 0 8 0 0 4096 0 23 0 0 17 2
217 88
188 88
0 0 9 0 0 8320 0 0 0 9 18 5
596 185
596 271
329 271
329 184
309 184
3 0 10 0 0 8320 0 6 0 0 26 3
463 31
463 19
188 19
0 1 9 0 0 0 0 0 2 10 0 2
584 185
600 185
2 2 9 0 0 0 0 1 4 0 0 4
568 169
584 169
584 200
568 200
3 3 11 0 0 4224 0 1 4 0 0 2
544 178
544 191
1 1 2 0 0 4096 0 4 3 0 0 2
544 227
544 241
1 1 2 0 0 4096 0 5 19 0 0 2
404 242
404 206
2 2 12 0 0 4224 0 19 6 0 0 3
404 170
404 51
451 51
2 1 5 0 0 4224 0 20 6 0 0 2
463 167
463 67
1 1 2 0 0 4096 0 7 20 0 0 2
463 241
463 203
1 3 8 0 0 4224 0 24 11 0 0 2
188 69
188 100
2 2 9 0 0 0 0 15 13 0 0 4
293 170
309 170
309 201
293 201
3 3 13 0 0 4224 0 15 13 0 0 2
269 179
269 192
1 1 2 0 0 0 0 13 14 0 0 2
269 228
269 242
1 1 2 0 0 0 0 12 22 0 0 2
129 243
129 207
2 2 14 0 0 4224 0 22 11 0 0 3
129 171
129 120
176 120
2 1 15 0 0 4224 0 21 11 0 0 2
188 168
188 136
1 1 2 0 0 0 0 10 21 0 0 2
188 242
188 204
1 2 2 0 0 4224 0 9 8 0 0 3
94 240
94 196
80 196
1 2 10 0 0 0 0 8 24 0 0 5
80 186
94 186
94 19
188 19
188 33
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.05 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

CircuitMaker Text
5.6
Probes: 1
U1A_1
Transient Analysis
0 279 195 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 110 10
176 83 1022 717
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 2 1
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 179 1190 496
9961490 0
0
6 Title:
5 Name:
0
0
0
32
9 Schottky~
219 22 55 0 2 5
0 6 5
0
0 0 848 90
6 1N6392
6 11 48 19
2 D1
15 -1 29 7
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 18
68 0 0 0 1 0 0 0
1 D
5130 0 0
2
5.89708e-315 0
0
9 Inductor~
219 133 111 0 2 5
0 6 3
0
0 0 848 0
5 430uH
-18 -17 17 -9
2 L1
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
391 0 0
2
42146 0
0
2 +V
167 334 141 0 1 3
0 8
0
0 0 53616 0
2 5V
-6 -13 8 -5
2 V7
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3124 0 0
2
42146 1
0
9 Schottky~
219 15 150 0 2 5
0 4 6
0
0 0 848 90
6 1N6392
12 -1 54 7
2 D2
26 -11 40 -3
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
3421 0 0
2
42146 2
0
10 Op-Amp5:A~
219 253 197 0 5 11
0 21 23 24 10 22
0
0 0 848 0
5 TL082
15 -25 50 -17
3 U1A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 3 0
1 U
8157 0 0
2
5.89708e-315 5.26354e-315
0
2 +V
167 253 225 0 1 3
0 10
0
0 0 53616 180
4 -15V
-13 -1 15 7
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5572 0 0
2
5.89708e-315 5.30499e-315
0
7 Ground~
168 419 315 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8901 0 0
2
5.89708e-315 5.32571e-315
0
2 +V
167 394 321 0 1 3
0 13
0
0 0 53616 180
4 -15V
-13 -1 15 7
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7361 0 0
2
5.89708e-315 5.34643e-315
0
9 2-In AND~
219 756 200 0 3 22
0 7 7 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
4747 0 0
2
5.89708e-315 5.3568e-315
0
2 +V
167 626 110 0 1 3
0 14
0
0 0 53616 0
2 5V
-6 -13 8 -5
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
972 0 0
2
5.89708e-315 5.36716e-315
0
2 +V
167 447 110 0 1 3
0 16
0
0 0 53616 0
2 5V
-6 -13 8 -5
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3472 0 0
2
5.89708e-315 5.37752e-315
0
12 NPN Trans:B~
219 842 200 0 3 7
0 18 19 2
0
0 0 848 0
6 BC547A
9 1 51 9
2 Q3
9 -11 23 -3
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
9998 0 0
2
5.89708e-315 5.38788e-315
0
7 Ground~
168 847 315 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3536 0 0
2
5.89708e-315 5.39306e-315
0
7 Ground~
168 615 315 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4597 0 0
2
5.89708e-315 5.39824e-315
0
5 4013~
219 660 227 0 6 22
0 2 14 17 11 9 7
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U3A
-12 -77 9 -69
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 0 2 1 1 0
1 U
3835 0 0
2
5.89708e-315 5.40342e-315
0
11 Signal Gen~
195 575 214 0 64 64
0 17 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1199715674 0 1084227584
0 814313567 814313567 930301191 930850946 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 66666.7 0 5 0 1e-09 1e-09 1.45e-05 1.5e-05 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
4 0/5V
-15 -30 13 -22
3 Osc
-10 -40 11 -32
0
0
42 %D %1 %2 DC 0 PULSE(0 5 0 1n 1n 14.5u 15u)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3670 0 0
2
5.89708e-315 5.4086e-315
0
2 +V
167 394 110 0 1 3
0 20
0
0 0 53616 0
3 15V
-9 -13 12 -5
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5616 0 0
2
5.89708e-315 5.41378e-315
0
12 Comparator6~
219 394 191 0 6 13
0 22 8 20 13 11 2
0
0 0 848 0
5 LM111
9 -19 44 -11
2 U2
8 -30 22 -22
0
0
23 %D %1 %2 %3 %4 %5 %6 %S
0
0
4 DIP8
13

0 2 3 8 4 7 1 2 3 8
4 7 1 0
88 0 0 256 1 0 0 0
1 U
9323 0 0
2
5.89708e-315 5.41896e-315
0
2 +V
167 253 110 0 1 3
0 24
0
0 0 53616 0
3 15V
-10 -13 11 -5
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
317 0 0
2
5.89708e-315 5.42414e-315
0
10 Capacitor~
219 127 229 0 2 5
0 2 21
0
0 0 848 90
5 100pF
10 0 45 8
2 C1
20 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3108 0 0
2
5.89708e-315 5.42933e-315
0
12 PNP Trans:B~
219 74 61 0 3 7
0 6 15 5
0
0 0 848 180
7 FZT790A
12 4 61 12
2 Q1
12 -12 26 -4
0
0
14 %D %1 %2 %3 %M
0
0
7 SOT-223
7

0 2 1 3 2 1 3 0
113 0 0 0 1 0 0 0
1 Q
4299 0 0
2
5.89708e-315 5.43192e-315
0
2 +V
167 63 17 0 1 3
0 5
0
0 0 53616 0
3 50V
-11 -14 10 -6
2 V0
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9672 0 0
2
5.89708e-315 5.43451e-315
0
7 Ground~
168 63 308 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7876 0 0
2
5.89708e-315 5.4371e-315
0
11 Resistor:A~
219 485 317 0 4 5
0 9 2 0 -1
0
0 0 880 270
3 10k
5 0 26 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6369 0 0
2
42146 3
0
9 Resistor~
219 128 163 0 2 5
0 3 4
0
0 0 880 180
4 0.68
-14 -14 14 -6
3 RS2
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9172 0 0
2
42146 4
0
11 Resistor:A~
219 803 200 0 2 5
0 12 19
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7100 0 0
2
5.89708e-315 5.43969e-315
0
11 Resistor:A~
219 847 154 0 2 5
0 18 15
0
0 0 880 602
2 1k
7 0 21 8
2 R7
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3820 0 0
2
5.89708e-315 5.44228e-315
0
11 Resistor:A~
219 182 260 0 4 5
0 23 2 0 -1
0
0 0 880 180
2 1k
-7 -15 7 -7
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7678 0 0
2
5.89708e-315 5.44487e-315
0
11 Resistor:A~
219 447 154 0 3 5
0 16 11 1
0
0 0 880 270
2 1k
8 0 22 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
961 0 0
2
5.89708e-315 5.44746e-315
0
11 Resistor:A~
219 249 260 0 2 5
0 23 22
0
0 0 880 0
2 9k
-7 -14 7 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3178 0 0
2
5.89708e-315 5.45005e-315
0
11 Resistor:A~
219 94 191 0 2 5
0 21 4
0
0 0 880 180
2 1k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3409 0 0
2
5.89708e-315 5.45264e-315
0
9 Resistor~
219 63 229 0 3 5
0 2 4 -1
0
0 0 880 90
3 0.1
5 0 26 8
3 RS1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3951 0 0
2
5.89708e-315 5.45523e-315
0
40
1 2 3 0 0 8320 0 25 2 0 0 4
146 163
175 163
175 111
151 111
2 1 4 0 0 8320 0 32 4 0 0 4
63 211
63 191
16 191
16 160
2 0 5 0 0 8320 0 1 0 0 11 5
23 42
23 30
62 30
62 31
63 31
1 1 6 0 0 8192 0 1 21 0 0 4
23 65
23 93
63 93
63 79
2 0 7 0 0 4096 0 9 0 0 18 3
732 209
713 209
713 191
1 0 6 0 0 4224 0 2 0 0 39 2
115 111
63 111
2 1 8 0 0 4224 0 18 3 0 0 3
376 185
334 185
334 150
1 5 9 0 0 8320 0 24 15 0 0 5
485 299
485 289
702 289
702 209
690 209
2 0 2 0 0 12288 0 24 0 0 15 5
485 335
485 348
446 348
446 294
419 294
2 0 4 0 0 0 0 25 0 0 38 3
110 163
63 163
63 191
1 3 5 0 0 0 0 22 21 0 0 2
63 26
63 43
4 1 10 0 0 0 0 5 6 0 0 2
253 210
253 210
1 0 2 0 0 4096 0 14 0 0 23 2
615 309
615 219
2 0 11 0 0 4096 0 29 0 0 19 2
447 172
447 183
1 6 2 0 0 4224 0 7 18 0 0 3
419 309
419 199
410 199
1 3 12 0 0 4224 0 26 9 0 0 2
785 200
777 200
1 4 13 0 0 4224 0 8 18 0 0 2
394 306
394 204
6 1 7 0 0 4224 0 15 9 0 0 2
684 191
732 191
5 4 11 0 0 12416 0 18 15 0 0 5
410 183
447 183
447 275
660 275
660 233
2 1 14 0 0 8320 0 15 10 0 0 3
636 191
626 191
626 119
2 2 15 0 0 8320 0 27 21 0 0 3
847 136
847 61
86 61
1 1 16 0 0 4224 0 11 29 0 0 2
447 119
447 136
1 2 2 0 0 0 0 15 16 0 0 5
660 170
660 163
615 163
615 219
606 219
1 3 17 0 0 4224 0 16 15 0 0 2
606 209
636 209
1 1 18 0 0 4224 0 12 27 0 0 2
847 182
847 172
1 3 2 0 0 0 0 13 12 0 0 2
847 309
847 218
2 2 19 0 0 4224 0 12 26 0 0 2
824 200
821 200
1 3 20 0 0 4224 0 17 18 0 0 2
394 119
394 178
1 0 2 0 0 0 0 20 0 0 30 2
127 238
127 260
2 0 2 0 0 0 0 28 0 0 40 2
164 260
63 260
1 0 21 0 0 4224 0 5 0 0 37 2
235 191
127 191
1 0 22 0 0 4224 0 18 0 0 34 2
376 197
279 197
1 0 23 0 0 4096 0 28 0 0 35 2
200 260
219 260
5 2 22 0 0 0 0 5 30 0 0 4
271 197
279 197
279 260
267 260
2 1 23 0 0 8320 0 5 30 0 0 4
235 203
219 203
219 260
231 260
1 3 24 0 0 4224 0 19 5 0 0 2
253 119
253 184
2 1 21 0 0 0 0 20 31 0 0 3
127 220
127 191
112 191
2 0 4 0 0 0 0 31 0 0 2 2
76 191
63 191
2 1 6 0 0 0 0 4 21 0 0 4
16 137
16 111
63 111
63 79
1 1 2 0 0 0 0 23 32 0 0 2
63 302
63 247
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 7.5e-05 3e-07 3e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

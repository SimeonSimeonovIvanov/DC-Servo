CircuitMaker Text
5.6
Probes: 1
U2_2
Transient Analysis
0 373 257 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 110 10
176 83 1022 717
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 2 1
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 179 457 276
9961490 0
0
6 Title:
5 Name:
0
0
0
39
11 Resistor:A~
219 163 130 0 4 5
0 7 2 0 -1
0
0 0 864 270
2 10
12 2 26 10
3 RL2
9 -11 30 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5130 0 0
2
42091.9 38
0
11 Resistor:A~
219 803 200 0 2 5
0 11 21
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
391 0 0
2
42091.9 37
0
11 Resistor:A~
219 847 154 0 2 5
0 20 17
0
0 0 864 602
2 1k
7 0 21 8
2 R7
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3124 0 0
2
42091.9 36
0
11 Resistor:A~
219 497 223 0 2 5
0 22 19
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3421 0 0
2
42091.9 35
0
11 Resistor:A~
219 182 260 0 4 5
0 9 2 0 -1
0
0 0 864 180
2 1k
-7 -15 7 -7
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8157 0 0
2
42091.9 34
0
11 Resistor:A~
219 447 154 0 3 5
0 18 3 1
0
0 0 864 270
2 1k
8 0 22 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5572 0 0
2
42091.9 33
0
11 Resistor:A~
219 249 260 0 2 5
0 9 8
0
0 0 864 0
2 9k
-7 -14 7 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8901 0 0
2
42091.9 32
0
11 Resistor:A~
219 94 191 0 2 5
0 24 6
0
0 0 864 180
2 1k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7361 0 0
2
42091.9 31
0
11 Resistor:A~
219 13 120 0 2 5
0 5 26
0
0 0 864 270
1 1
17 3 24 11
3 RL1
10 -9 31 -1
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4747 0 0
2
42091.9 30
0
9 Resistor~
219 63 229 0 3 5
0 2 6 -1
0
0 0 864 90
3 0.1
5 0 26 8
3 RS1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
972 0 0
2
42091.9 29
0
12 Transformer~
219 88 135 0 4 9
0 7 2 5 6
0
0 0 576 512
0
2 T1
-7 -30 7 -22
0
0
49 LP%D %1 %2 2mh
LS%D %3 %4 2mh
%D LP%D LS%D .999
0
0
0
9

0 1 2 3 4 1 2 3 4 0
75 0 0 0 1 0 0 0
1 T
3472 0 0
2
42091.9 28
0
7 Ground~
168 138 173 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9998 0 0
2
42091.9 27
0
10 Capacitor~
219 250 299 0 2 5
0 8 9
0
0 0 832 180
5 330pF
-16 -18 19 -10
2 C2
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3536 0 0
2
42091.9 26
0
10 Op-Amp5:A~
219 253 197 0 5 11
0 24 9 25 10 8
0
0 0 832 0
5 TL082
15 -25 50 -17
3 U1A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 3 0
1 U
4597 0 0
2
42091.9 25
0
2 +V
167 253 225 0 1 3
0 10
0
0 0 53600 180
4 -15V
-13 -1 15 7
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3835 0 0
2
42091.9 24
0
7 Ground~
168 447 315 0 1 3
0 2
0
0 0 53344 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3670 0 0
2
42091.9 23
0
7 Ground~
168 419 315 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5616 0 0
2
42091.9 22
0
2 +V
167 394 321 0 1 3
0 12
0
0 0 53600 180
4 -15V
-13 -1 15 7
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9323 0 0
2
42091.9 21
0
9 2-In AND~
219 756 200 0 3 22
0 13 14 11
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
317 0 0
2
42091.9 20
0
2 +V
167 626 110 0 1 3
0 16
0
0 0 53600 0
2 5V
-6 -13 8 -5
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3108 0 0
2
42091.9 19
0
2 +V
167 447 110 0 1 3
0 18
0
0 0 53600 0
2 5V
-6 -13 8 -5
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4299 0 0
2
42091.9 18
0
12 NPN Trans:B~
219 842 200 0 3 7
0 20 21 2
0
0 0 832 0
6 BC547A
9 1 51 9
2 Q3
9 -11 23 -3
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
9672 0 0
2
42091.9 17
0
7 Ground~
168 847 315 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7876 0 0
2
42091.9 16
0
7 Ground~
168 615 315 0 1 3
0 2
0
0 0 53344 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6369 0 0
2
42091.9 15
0
5 4013~
219 660 227 0 6 22
0 2 16 14 3 19 13
0
0 0 4704 0
4 4013
10 -60 38 -52
3 U3A
-12 -77 9 -69
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 0 2 1 1 0
1 U
9172 0 0
2
42091.9 14
0
11 Signal Gen~
195 575 214 0 64 64
0 14 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1176256512 0 1084227584
0 814313567 814313567 952580797 953267991 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 10000 0 5 0 1e-09 1e-09 9.5e-05 0.0001 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
4 0/5V
-15 -30 13 -22
3 Osc
-10 -40 11 -32
0
0
41 %D %1 %2 DC 0 PULSE(0 5 0 1n 1n 95u 100u)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
7100 0 0
2
42091.9 13
0
12 NPN Trans:B~
219 456 223 0 3 7
0 3 22 2
0
0 0 832 512
6 BC547A
-2 14 40 22
2 Q2
6 -10 20 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
3820 0 0
2
42091.9 12
0
2 +V
167 311 187 0 1 3
0 2
0
0 0 54112 90
4 2.5V
-10 -17 18 -9
4 Ref1
-10 -29 18 -21
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7678 0 0
2
42091.9 11
0
11 Signal Gen~
195 315 255 0 64 64
0 15 2 2 86 -9 9 0 0 0
0 0 0 0 0 0 0 1120403456 1075838976 1075838976
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 100 2.5 2.5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
4 0/5V
-15 -30 13 -22
3 Ref
-10 -40 11 -32
0
0
34 %D %1 %2 DC 0 SIN(2.5 2.5 100 0 0)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
961 0 0
2
42091.9 10
0
7 Ground~
168 354 315 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3178 0 0
2
42091.9 9
0
2 +V
167 394 110 0 1 3
0 23
0
0 0 53600 0
3 15V
-9 -13 12 -5
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3409 0 0
2
42091.9 8
0
12 Comparator6~
219 394 191 0 6 13
0 8 15 23 12 3 2
0
0 0 832 0
5 LM111
9 -19 44 -11
2 U2
8 -30 22 -22
0
0
23 %D %1 %2 %3 %4 %5 %6 %S
0
0
4 DIP8
13

0 2 3 8 4 7 1 2 3 8
4 7 1 0
88 0 0 256 1 0 0 0
1 U
3951 0 0
2
42091.9 7
0
2 +V
167 253 110 0 1 3
0 25
0
0 0 53600 0
3 15V
-10 -13 11 -5
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8885 0 0
2
42091.9 6
0
10 Capacitor~
219 127 229 0 2 5
0 2 24
0
0 0 832 90
5 100nF
12 0 47 8
2 C1
20 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3780 0 0
2
42091.9 5
0
10 Capacitor~
219 13 162 0 2 5
0 6 26
0
0 0 832 90
4 10nF
14 3 42 11
3 CL1
15 -7 36 1
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9265 0 0
2
42091.9 4
0
9 Schottky~
219 12 62 0 2 5
0 5 4
0
0 0 832 90
6 1N5828
6 11 48 19
2 D1
15 -1 29 7
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
9442 0 0
2
42091.9 3
0
12 PNP Trans:B~
219 74 61 0 3 7
0 5 17 4
0
0 0 832 180
7 FZT790A
12 4 61 12
2 Q1
12 -12 26 -4
0
0
14 %D %1 %2 %3 %M
0
0
7 SOT-223
7

0 2 1 3 2 1 3 0
113 0 0 0 1 0 0 0
1 Q
9424 0 0
2
42091.9 2
0
2 +V
167 63 17 0 1 3
0 4
0
0 0 53600 0
3 36V
-11 -14 10 -6
2 V0
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9968 0 0
2
42091.9 1
0
7 Ground~
168 63 308 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9281 0 0
2
42091.9 0
0
49
1 0 3 0 0 16 0 27 0 0 14 2
447 205
447 183
2 0 4 0 0 16 0 36 0 0 3 3
13 49
13 34
63 34
1 3 4 0 0 16 0 38 37 0 0 2
63 26
63 43
1 0 5 0 0 16 0 36 0 0 48 2
13 72
13 91
1 0 2 0 0 16 0 12 0 0 8 2
138 167
138 162
4 0 6 0 0 16 0 11 0 0 45 3
69 151
63 151
63 191
3 0 5 0 0 16 0 11 0 0 48 3
69 119
63 119
63 89
2 2 2 0 0 16 0 1 11 0 0 5
163 148
163 162
114 162
114 143
107 143
1 1 7 0 0 16 0 1 11 0 0 5
163 112
163 99
113 99
113 127
107 127
1 0 8 0 0 16 0 13 0 0 41 3
259 299
279 299
279 260
2 0 9 0 0 16 0 13 0 0 40 3
241 299
219 299
219 260
4 1 10 0 0 16 0 14 15 0 0 2
253 210
253 210
1 0 2 0 0 16 0 24 0 0 29 2
615 309
615 219
2 0 3 0 0 16 0 6 0 0 23 2
447 172
447 183
1 3 2 0 0 16 0 16 27 0 0 2
447 309
447 241
1 6 2 0 0 16 0 17 32 0 0 3
419 309
419 199
410 199
1 3 11 0 0 16 0 2 19 0 0 2
785 200
777 200
1 4 12 0 0 16 0 18 32 0 0 2
394 306
394 204
1 0 2 0 0 16 0 30 0 0 21 2
354 309
354 260
6 1 13 0 0 16 0 25 19 0 0 2
684 191
732 191
1 2 2 0 0 16 0 28 29 0 0 4
322 185
354 185
354 260
346 260
2 0 14 0 0 16 0 19 0 0 30 5
732 209
715 209
715 302
626 302
626 209
5 4 3 0 0 16 0 32 25 0 0 5
410 183
538 183
538 279
660 279
660 233
1 2 15 0 0 16 0 29 32 0 0 4
346 250
364 250
364 185
376 185
2 1 16 0 0 16 0 25 20 0 0 3
636 191
626 191
626 119
2 2 17 0 0 16 0 3 37 0 0 3
847 136
847 61
86 61
1 1 18 0 0 16 0 21 6 0 0 2
447 119
447 136
2 5 19 0 0 16 0 4 25 0 0 6
515 223
527 223
527 290
700 290
700 209
690 209
1 2 2 0 0 16 0 25 26 0 0 5
660 170
660 163
615 163
615 219
606 219
1 3 14 0 0 16 0 26 25 0 0 2
606 209
636 209
1 1 20 0 0 16 0 22 3 0 0 2
847 182
847 172
1 3 2 0 0 16 0 23 22 0 0 2
847 309
847 218
2 2 21 0 0 16 0 22 2 0 0 2
824 200
821 200
1 2 22 0 0 16 0 4 27 0 0 2
479 223
470 223
1 3 23 0 0 16 0 31 32 0 0 2
394 119
394 178
1 0 2 0 0 16 0 34 0 0 37 2
127 238
127 260
2 0 2 0 0 16 0 5 0 0 49 2
164 260
63 260
1 0 24 0 0 16 0 14 0 0 44 2
235 191
127 191
1 0 8 0 0 16 0 32 0 0 41 2
376 197
279 197
1 0 9 0 0 16 0 5 0 0 42 2
200 260
219 260
5 2 8 0 0 16 0 14 7 0 0 4
271 197
279 197
279 260
267 260
2 1 9 0 0 16 0 14 7 0 0 4
235 203
219 203
219 260
231 260
1 3 25 0 0 16 0 33 14 0 0 2
253 119
253 184
2 1 24 0 0 16 0 34 8 0 0 3
127 220
127 191
112 191
2 0 6 0 0 16 0 8 0 0 47 2
76 191
63 191
2 2 26 0 0 16 0 35 9 0 0 2
13 153
13 138
1 2 6 0 0 16 0 35 10 0 0 4
13 171
13 191
63 191
63 211
1 1 5 0 0 16 0 9 37 0 0 4
13 102
13 90
63 90
63 79
1 1 2 0 0 16 0 39 10 0 0 2
63 302
63 247
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.05 5e-05 5e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

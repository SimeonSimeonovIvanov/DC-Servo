CircuitMaker Text
5.6
Probes: 1
R1_2
Operating Point
0 385 116 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 31 14 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 170 10
176 83 1022 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 2 0
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 179 457 276
9961490 0
0
2 

2 

0
0
0
4
9 V Source~
197 77 110 0 2 5
0 3 2
0
0 0 18016 0
3 10V
13 0 34 8
7 Voltage
-64 -12 -15 -4
6 Source
-61 2 -19 10
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
6118 0 0
2
42092.2 3
0
9 V Source~
197 260 158 0 2 5
0 5 2
0
0 0 17632 0
3 10V
13 0 34 8
3 Vs2
13 -10 34 -2
8 Back EMF
19 -3 75 5
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
34 0 0
2
42092.2 2
0
8 Coil 3T~
219 260 110 0 2 5
0 4 5
0
0 0 1088 270
3 1uH
8 -1 29 7
2 L1
12 -11 26 -3
1 L
13 -3 20 5
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
6357 0 0
2
42092.2 1
0
11 Resistor:A~
219 260 63 0 2 5
0 3 4
0
0 0 1120 270
2 1k
8 0 22 8
2 R1
8 -10 22 -2
1 R
13 -4 20 4
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
319 0 0
2
42092.2 0
0
4
2 2 2 0 0 16 0 2 1 0 0 4
260 179
260 188
77 188
77 131
1 1 3 0 0 16 0 4 1 0 0 4
260 45
260 37
77 37
77 89
2 1 4 0 0 16 0 4 3 0 0 2
260 81
260 90
2 1 5 0 0 16 0 3 2 0 0 2
260 130
260 137
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
110 8 236 32
112 11 233 27
15 M = Km * I [Nm]
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
100 99 251 123
103 102 247 118
18 P = Speed * Tm [W]
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
206 198 333 222
209 201 329 217
15 Vb = Kb * Speed
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
7 198 157 219
10 202 153 217
17 Vs = Vr + Vl + Vb
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
292 53 377 77
294 55 374 71
10 Vr = I * R
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
296 101 461 125
298 103 458 119
20 Vl = L * ( dI / dt )
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

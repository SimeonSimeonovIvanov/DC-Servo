CircuitMaker Text
5.6
Probes: 1
U1A_1
Transient Analysis
0 307 200 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 130 10
176 79 1918 1019
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 2 1
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 2086 645
9961490 0
0
6 Title:
5 Name:
0
0
0
38
10 Capacitor~
219 249 303 0 2 5
0 4 5
0
0 0 848 180
5 330pF
-16 -18 19 -10
2 C3
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7519 0 0
2
5.89662e-315 0
0
10 Op-Amp5:A~
219 252 201 0 5 11
0 20 5 21 6 4
0
0 0 848 0
5 TL082
15 -25 50 -17
3 U1A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 3 0
1 U
377 0 0
2
5.89662e-315 0
0
2 +V
167 252 229 0 1 3
0 6
0
0 0 53616 180
4 -15V
-13 -1 15 7
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8816 0 0
2
5.89662e-315 0
0
7 Ground~
168 446 319 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3877 0 0
2
5.89662e-315 0
0
7 Ground~
168 418 319 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
926 0 0
2
5.89662e-315 0
0
2 +V
167 393 325 0 1 3
0 8
0
0 0 53616 180
4 -15V
-13 -1 15 7
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7262 0 0
2
5.89662e-315 0
0
9 2-In AND~
219 738 204 0 3 22
0 9 10 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
5267 0 0
2
43873.9 0
0
10 Capacitor~
219 186 303 0 2 5
0 2 2
0
0 0 848 180
3 1pF
-10 -18 11 -10
2 C2
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
8838 0 0
2
43873.9 1
0
2 +V
167 625 114 0 1 3
0 12
0
0 0 53616 0
2 5V
-6 -13 8 -5
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7159 0 0
2
43873.9 2
0
2 +V
167 446 114 0 1 3
0 14
0
0 0 53616 0
2 5V
-6 -13 8 -5
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5812 0 0
2
43873.9 3
0
12 NPN Trans:B~
219 841 204 0 3 7
0 16 17 2
0
0 0 848 0
6 BC547A
9 1 51 9
2 Q3
9 -11 23 -3
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
331 0 0
2
43873.9 4
0
7 Ground~
168 846 319 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9604 0 0
2
43873.9 5
0
7 Ground~
168 614 319 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7518 0 0
2
43873.9 6
0
5 4013~
219 659 231 0 6 22
0 2 12 10 3 15 9
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U3A
-12 -77 9 -69
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 0 2 1 1 0
1 U
4832 0 0
2
43873.9 7
0
11 Signal Gen~
195 574 218 0 64 64
0 10 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1176256512 0 1084227584
0 814313567 814313567 952580797 953267991 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 10000 0 5 0 1e-09 1e-09 9.5e-05 0.0001 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
4 0/5V
-15 -30 13 -22
3 Osc
-10 -40 11 -32
0
0
41 %D %1 %2 DC 0 PULSE(0 5 0 1n 1n 95u 100u)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
6798 0 0
2
43873.9 8
0
12 NPN Trans:B~
219 455 227 0 3 7
0 3 18 2
0
0 0 848 512
6 BC547A
-2 14 40 22
2 Q2
6 -10 20 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
3336 0 0
2
43873.9 9
0
2 +V
167 310 191 0 1 3
0 2
0
0 0 54128 90
4 2.5V
-10 -17 18 -9
4 Ref1
-10 -29 18 -21
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8370 0 0
2
43873.9 10
0
11 Signal Gen~
195 314 259 0 64 64
0 11 2 2 86 -9 9 0 0 0
0 0 0 0 0 0 0 1120403456 1075838976 1075838976
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 100 2.5 2.5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
4 0/5V
-15 -30 13 -22
3 Ref
-10 -40 11 -32
0
0
34 %D %1 %2 DC 0 SIN(2.5 2.5 100 0 0)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3910 0 0
2
43873.9 11
0
7 Ground~
168 353 319 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
316 0 0
2
43873.9 12
0
2 +V
167 393 114 0 1 3
0 19
0
0 0 53616 0
3 15V
-9 -13 12 -5
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
536 0 0
2
43873.9 13
0
12 Comparator6~
219 393 195 0 6 13
0 4 11 19 8 3 2
0
0 0 848 0
5 LM111
9 -19 44 -11
2 U2
8 -30 22 -22
0
0
23 %D %1 %2 %3 %4 %5 %6 %S
0
0
4 DIP8
13

0 2 3 8 4 7 1 2 3 8
4 7 1 0
88 0 0 256 1 0 0 0
1 U
4460 0 0
2
43873.9 14
0
2 +V
167 252 114 0 1 3
0 21
0
0 0 53616 0
3 15V
-10 -13 11 -5
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3260 0 0
2
43873.9 15
0
10 Capacitor~
219 126 233 0 2 5
0 2 20
0
0 0 848 90
5 4.7nF
12 0 47 8
2 C1
20 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5156 0 0
2
43873.9 16
0
10 Capacitor~
219 12 166 0 2 5
0 22 24
0
0 0 848 90
4 47nF
13 0 41 8
3 CL1
12 -10 33 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3133 0 0
2
43873.9 17
0
8 Coil 3T~
219 62 144 0 2 5
0 23 22
0
0 0 848 782
3 1mH
8 0 29 8
2 L1
9 -10 23 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
5523 0 0
2
5.89662e-315 0
0
9 Schottky~
219 11 66 0 2 5
0 23 25
0
0 0 848 90
6 1N5828
6 7 48 15
2 D1
6 -16 20 -8
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
3746 0 0
2
5.89662e-315 5.26354e-315
0
12 PNP Trans:B~
219 73 65 0 3 7
0 23 13 25
0
0 0 848 180
7 FZT790A
12 4 61 12
2 Q1
12 -12 26 -4
0
0
14 %D %1 %2 %3 %M
0
0
7 SOT-223
7

0 2 1 3 2 1 3 0
113 0 0 0 1 0 0 0
1 Q
5668 0 0
2
5.89662e-315 5.30499e-315
0
2 +V
167 62 17 0 1 3
0 25
0
0 0 53616 0
3 36V
-11 -14 10 -6
2 V0
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5368 0 0
2
5.89662e-315 5.32571e-315
0
7 Ground~
168 62 312 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8293 0 0
2
5.89662e-315 5.34643e-315
0
11 Resistor:A~
219 802 204 0 2 5
0 7 17
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3232 0 0
2
43873.9 18
0
11 Resistor:A~
219 846 158 0 2 5
0 16 13
0
0 0 880 602
2 1k
7 0 21 8
2 R7
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6644 0 0
2
43873.9 19
0
11 Resistor:A~
219 496 227 0 2 5
0 18 15
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4978 0 0
2
43873.9 20
0
11 Resistor:A~
219 181 264 0 4 5
0 5 2 0 -1
0
0 0 880 180
2 1k
-7 -15 7 -7
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9207 0 0
2
43873.9 21
0
11 Resistor:A~
219 446 158 0 3 5
0 14 3 1
0
0 0 880 270
2 1k
8 0 22 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6998 0 0
2
43873.9 22
0
11 Resistor:A~
219 248 264 0 2 5
0 5 4
0
0 0 880 0
2 9k
-7 -14 7 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3175 0 0
2
43873.9 23
0
11 Resistor:A~
219 93 195 0 2 5
0 20 22
0
0 0 880 180
2 1k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3378 0 0
2
43873.9 24
0
11 Resistor:A~
219 12 124 0 2 5
0 23 24
0
0 0 880 270
3 0.5
5 0 26 8
3 RL1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
922 0 0
2
43873.9 25
0
9 Resistor~
219 62 233 0 3 5
0 2 22 -1
0
0 0 880 90
3 0.1
5 0 26 8
3 RS1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6891 0 0
2
5.89662e-315 5.3568e-315
0
48
1 0 3 0 0 4096 0 16 0 0 6 2
446 209
446 188
1 0 4 0 0 8192 0 1 0 0 35 3
258 303
278 303
278 264
2 0 5 0 0 8192 0 1 0 0 34 3
240 303
218 303
218 264
4 1 6 0 0 0 0 2 3 0 0 2
252 214
252 214
1 0 2 0 0 4096 0 13 0 0 23 2
614 313
614 223
2 0 3 0 0 0 0 34 0 0 16 2
446 176
446 187
1 3 2 0 0 0 0 4 16 0 0 2
446 313
446 245
1 6 2 0 0 4224 0 5 21 0 0 3
418 313
418 203
409 203
1 3 7 0 0 4224 0 30 7 0 0 2
784 204
759 204
1 4 8 0 0 4224 0 6 21 0 0 2
393 310
393 208
1 0 2 0 0 0 0 19 0 0 14 2
353 313
353 264
1 0 2 0 0 0 0 8 0 0 18 5
195 303
206 303
206 324
126 324
126 303
6 1 9 0 0 4224 0 14 7 0 0 2
683 195
714 195
1 2 2 0 0 0 0 17 18 0 0 4
321 189
353 189
353 264
345 264
2 0 10 0 0 8320 0 7 0 0 24 5
714 213
707 213
707 306
625 306
625 213
5 4 3 0 0 4224 0 21 14 0 0 5
409 187
537 187
537 283
659 283
659 237
1 2 11 0 0 8320 0 18 21 0 0 4
345 254
363 254
363 189
375 189
2 0 2 0 0 0 0 8 0 0 30 3
177 303
126 303
126 264
2 1 12 0 0 8320 0 14 9 0 0 3
635 195
625 195
625 123
2 2 13 0 0 8320 0 31 27 0 0 3
846 140
846 65
85 65
1 1 14 0 0 4224 0 10 34 0 0 2
446 123
446 140
2 5 15 0 0 12416 0 32 14 0 0 6
514 227
526 227
526 294
696 294
696 213
689 213
1 2 2 0 0 0 0 14 15 0 0 5
659 174
659 167
614 167
614 223
605 223
1 3 10 0 0 0 0 15 14 0 0 2
605 213
635 213
1 1 16 0 0 4224 0 11 31 0 0 2
846 186
846 176
1 3 2 0 0 0 0 12 11 0 0 2
846 313
846 222
2 2 17 0 0 4224 0 11 30 0 0 2
823 204
820 204
1 2 18 0 0 4224 0 32 16 0 0 2
478 227
469 227
1 3 19 0 0 4224 0 20 21 0 0 2
393 123
393 182
1 0 2 0 0 0 0 23 0 0 31 2
126 242
126 264
2 0 2 0 0 0 0 33 0 0 48 2
163 264
62 264
1 0 20 0 0 4224 0 2 0 0 38 2
234 195
126 195
1 0 4 0 0 4224 0 21 0 0 35 2
375 201
278 201
1 0 5 0 0 0 0 33 0 0 36 2
199 264
218 264
5 2 4 0 0 0 0 2 35 0 0 4
270 201
278 201
278 264
266 264
2 1 5 0 0 8320 0 2 35 0 0 4
234 207
218 207
218 264
230 264
1 3 21 0 0 4224 0 22 2 0 0 2
252 123
252 188
2 1 20 0 0 0 0 23 36 0 0 3
126 224
126 195
111 195
2 0 22 0 0 4096 0 36 0 0 41 2
75 195
62 195
1 0 23 0 0 4096 0 37 0 0 44 2
12 106
12 94
1 0 22 0 0 8192 0 24 0 0 43 3
12 175
12 195
62 195
2 2 24 0 0 4224 0 24 37 0 0 2
12 157
12 142
2 2 22 0 0 4224 0 38 25 0 0 2
62 215
62 164
1 0 23 0 0 8320 0 26 0 0 46 3
12 76
12 94
62 94
2 0 25 0 0 8320 0 26 0 0 47 3
12 53
12 37
62 37
1 1 23 0 0 0 0 25 27 0 0 2
62 124
62 83
1 3 25 0 0 0 0 28 27 0 0 2
62 26
62 47
1 1 2 0 0 0 0 29 38 0 0 2
62 306
62 251
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.02 0.0001 0.0001
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

CircuitMaker Text
5.6
Probes: 1
U2_5
Transient Analysis
0 321 78 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 200 10
176 83 1022 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 2 1
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 179 1190 496
9961490 0
0
6 Title:
5 Name:
0
0
0
18
7 Ground~
168 110 211 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3978 0 0
2
42166 13
0
8 Op-Amp5~
219 137 138 0 5 11
0 7 6 9 8 5
0
0 0 848 0
5 TL082
15 -25 50 -17
3 U1A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 0 2 1 1 0
1 U
3494 0 0
2
42166 12
0
2 +V
167 137 166 0 1 3
0 8
0
0 0 53616 180
4 -15V
-14 0 14 8
2 V9
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3507 0 0
2
42166 11
0
2 +V
167 137 116 0 1 3
0 9
0
0 0 53616 0
4 +15V
-13 -14 15 -6
2 V8
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5151 0 0
2
42166 10
0
12 Comparator6~
219 269 98 0 6 13
0 3 4 13 11 15 16
0
0 0 848 0
5 LM111
15 -25 50 -17
2 U2
26 -35 40 -27
0
0
23 %D %1 %2 %3 %4 %5 %6 %S
0
0
0
13

0 1 2 3 4 5 6 1 2 3
4 5 6 0
88 0 0 0 1 0 0 0
1 U
3701 0 0
2
42166 9
0
12 Comparator6~
219 269 180 0 6 13
0 5 3 14 12 16 2
0
0 0 848 0
5 LM111
15 -25 50 -17
2 U3
26 -35 40 -27
0
0
23 %D %1 %2 %3 %4 %5 %6 %S
0
0
0
13

0 1 2 3 4 5 6 1 2 3
4 5 6 0
88 0 0 0 1 0 0 0
1 U
8585 0 0
2
42166 8
0
2 +V
167 269 158 0 1 3
0 14
0
0 0 53616 0
4 +15V
-13 -14 15 -6
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8809 0 0
2
42166 7
0
2 +V
167 269 76 0 1 3
0 13
0
0 0 53616 0
4 +15V
-13 -14 15 -6
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5993 0 0
2
42166 6
0
2 +V
167 269 208 0 1 3
0 12
0
0 0 53616 180
4 -15V
-14 0 14 8
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8654 0 0
2
42166 5
0
2 +V
167 269 126 0 1 3
0 11
0
0 0 53616 180
4 -15V
-14 0 14 8
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7223 0 0
2
42166 4
0
7 Ground~
168 321 211 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3641 0 0
2
42166 3
0
2 +V
167 321 17 0 1 3
0 10
0
0 0 53616 0
3 +5V
-10 -15 11 -7
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3104 0 0
2
42166 2
0
2 +V
167 213 140 0 1 3
0 3
0
0 0 54128 90
2 3V
-6 5 8 13
2 FB
-5 -16 9 -8
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3296 0 0
2
42166 1
0
2 +V
167 26 134 0 1 3
0 4
0
0 0 55152 90
4 3.5V
-11 7 17 15
2 SP
-5 -17 9 -9
8 SP >= 0V
-24 22 32 30
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8534 0 0
2
42166 0
0
11 Resistor:A~
219 110 179 0 4 5
0 7 2 0 -1
0
0 0 880 270
4 5.1k
-35 -2 -7 6
2 R3
-28 -13 -14 -5
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
949 0 0
2
42166 17
0
11 Resistor:A~
219 138 92 0 2 5
0 5 6
0
0 0 880 180
3 10k
-11 -14 10 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3371 0 0
2
42166 16
0
11 Resistor:A~
219 82 132 0 4 5
0 6 4 0 1
0
0 0 880 180
3 10k
-11 -14 10 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7311 0 0
2
42166 15
0
11 Resistor:A~
219 321 55 0 4 5
0 15 10 0 1
0
0 0 880 90
4 5.1k
10 1 38 9
2 R4
16 -10 30 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3409 0 0
2
42166 14
0
20
2 0 3 0 0 8336 0 6 0 0 3 3
251 174
239 174
239 138
2 0 4 0 0 12432 0 5 0 0 4 5
251 92
239 92
239 62
51 62
51 132
1 1 3 0 0 16 0 5 13 0 0 4
251 104
239 104
239 138
224 138
1 2 4 0 0 16 0 14 17 0 0 2
37 132
64 132
0 1 5 0 0 8336 0 0 6 6 0 3
188 138
188 186
251 186
1 5 5 0 0 16 0 16 2 0 0 4
156 92
188 92
188 138
155 138
2 1 2 0 0 4112 0 15 1 0 0 2
110 197
110 205
2 0 6 0 0 8336 0 16 0 0 12 3
120 92
110 92
110 132
1 1 7 0 0 4240 0 15 2 0 0 3
110 161
110 144
119 144
1 4 8 0 0 16 0 3 2 0 0 2
137 151
137 151
1 3 9 0 0 16 0 4 2 0 0 2
137 125
137 125
1 2 6 0 0 16 0 17 2 0 0 2
100 132
119 132
1 2 10 0 0 4240 0 12 18 0 0 2
321 26
321 37
1 6 2 0 0 8336 0 11 6 0 0 3
321 205
321 188
285 188
1 4 11 0 0 16 0 10 5 0 0 2
269 111
269 111
1 4 12 0 0 16 0 9 6 0 0 2
269 193
269 193
1 3 13 0 0 16 0 8 5 0 0 2
269 85
269 85
1 3 14 0 0 16 0 7 6 0 0 2
269 167
269 167
1 5 15 0 0 8336 0 18 5 0 0 3
321 73
321 90
285 90
6 5 16 0 0 8336 0 5 6 0 0 4
285 106
321 106
321 172
285 172
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 240 10
176 83 1022 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 2 0
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
5 4 0.309148 0.500000
344 179 457 276
42991634 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 14 154 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 PWM
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7168 0 0
2
5.89666e-315 5.30499e-315
0
13 Logic Switch~
5 206 229 0 1 11
0 7
0
0 0 21360 90
2 0V
11 0 25 8
2 V1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3171 0 0
2
5.89666e-315 5.26354e-315
0
13 Logic Switch~
5 14 99 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 FB
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4139 0 0
2
5.89666e-315 0
0
14 Logic Display~
6 251 75 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 G3L
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6435 0 0
2
5.89666e-315 5.39306e-315
0
14 Logic Display~
6 316 74 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 G4L
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5283 0 0
2
5.89666e-315 5.38788e-315
0
9 Inverter~
13 65 189 0 2 22
0 8 6
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
6874 0 0
2
5.89666e-315 5.37752e-315
0
5 4013~
219 147 225 0 6 22
0 7 6 9 8 2 3
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U1B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 0 2 2 1 0
1 U
5305 0 0
2
5.89666e-315 5.36716e-315
0
5 4013~
219 147 135 0 6 22
0 7 8 9 6 4 5
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U1A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 0 2 1 1 0
1 U
34 0 0
2
5.89666e-315 5.3568e-315
0
14 Logic Display~
6 251 23 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 G1H
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
969 0 0
2
5.89666e-315 5.34643e-315
0
14 Logic Display~
6 316 23 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 G2H
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8402 0 0
2
5.89666e-315 5.32571e-315
0
13
5 1 2 0 0 4224 0 7 10 0 0 5
177 207
339 207
339 47
316 47
316 41
6 1 3 0 0 8320 0 7 4 0 0 3
171 189
251 189
251 93
5 1 4 0 0 8320 0 8 9 0 0 5
177 117
228 117
228 47
251 47
251 41
6 1 5 0 0 4224 0 8 5 0 0 3
171 99
316 99
316 92
4 0 6 0 0 12432 0 8 0 0 13 4
147 141
147 145
113 145
113 189
1 0 7 0 0 4096 0 2 0 0 8 2
207 216
207 158
4 0 8 0 0 8320 0 7 0 0 12 4
147 231
147 241
39 241
39 189
1 1 7 0 0 12416 0 7 8 0 0 6
147 168
147 158
207 158
207 68
147 68
147 78
1 0 9 0 0 4096 0 1 0 0 11 2
26 154
100 154
1 0 8 0 0 0 0 3 0 0 12 2
26 99
39 99
3 3 9 0 0 8320 0 8 7 0 0 4
123 117
100 117
100 207
123 207
2 1 8 0 0 0 0 8 6 0 0 4
123 99
39 99
39 189
50 189
2 2 6 0 0 0 0 6 7 0 0 6
86 189
113 189
113 187
113 187
113 189
123 189
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

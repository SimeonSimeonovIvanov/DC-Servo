CircuitMaker Text
5.6
Probes: 1
C2_2
Transient Analysis
0 308 176 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 130 10
176 83 1022 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 2 0
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 179 1190 496
9961490 0
0
6 Title:
5 Name:
0
0
0
39
10 Capacitor~
219 274 32 0 2 5
0 6 5
0
0 0 848 0
5 0.1nF
-18 -18 17 -10
2 C2
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7128 0 0
2
41826.7 0
0
10 Capacitor~
219 277 110 0 2 5
0 4 3
0
0 0 848 0
5 220nF
-18 -18 17 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5367 0 0
2
41826.7 1
0
7 Ground~
168 145 193 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7140 0 0
2
41826.7 2
0
7 Ground~
168 190 193 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4903 0 0
2
41826.7 3
0
8 Op-Amp5~
219 216 172 0 5 11
0 2 6 25 24 10
0
0 0 848 0
5 TL082
-39 -28 -4 -20
3 U2A
-33 -39 -12 -31
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 2 0
1 U
3690 0 0
2
41826.7 4
0
2 +V
167 216 136 0 1 3
0 25
0
0 0 53616 0
4 +15V
-14 -14 14 -6
2 V7
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8598 0 0
2
41826.7 5
0
2 +V
167 216 213 0 1 3
0 24
0
0 0 53616 180
4 -15V
-12 -1 16 7
2 V6
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5737 0 0
2
41826.7 6
0
11 Signal Gen~
195 86 171 0 64 64
0 23 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1101004800 -1119040307 1028443341
0 814313567 814313567 1020054733 1028443341 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 20 -0.05 0.05 0 1e-09 1e-09 0.025 0.05 0
0 0 0 0 0 0 0 0 0 0
0
0 0 1360 0
9 -50m/50mV
-33 -30 30 -22
2 V5
-7 -40 7 -32
8 Speed SP
-27 -40 29 -32
0
45 %D %1 %2 DC 0 PULSE(-50m 50m 0 1n 1n 25m 50m)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3882 0 0
2
41826.7 7
0
2 +V
167 26 362 0 1 3
0 11
0
0 0 53616 90
2 6V
-7 -15 7 -7
2 V8
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3440 0 0
2
41826.7 8
0
2 +V
167 282 394 0 1 3
0 21
0
0 0 53616 180
4 -15V
-12 -1 16 7
2 V3
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5176 0 0
2
41826.7 9
0
2 +V
167 282 342 0 1 3
0 22
0
0 0 53616 0
4 +15V
-14 -14 14 -6
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9582 0 0
2
41826.7 10
0
8 Op-Amp5~
219 282 365 0 5 11
0 20 18 22 21 19
0
0 0 848 0
5 TL082
15 -25 50 -17
3 U2B
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 5 6 8 4 7 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 2 2 0
1 U
9862 0 0
2
41826.7 11
0
7 Ground~
168 256 466 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5432 0 0
2
41826.7 12
0
7 Ground~
168 335 466 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3602 0 0
2
41826.7 13
0
7 Ground~
168 165 466 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4714 0 0
2
41826.7 14
0
2 +V
167 112 395 0 1 3
0 16
0
0 0 53616 180
4 -15V
-12 -1 16 7
2 V2
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3834 0 0
2
41826.7 15
0
2 +V
167 112 343 0 1 3
0 17
0
0 0 53616 0
4 +15V
-14 -14 14 -6
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3577 0 0
2
41826.7 16
0
8 Op-Amp5~
219 112 366 0 5 11
0 14 15 17 16 12
0
0 0 848 0
5 TL082
15 -25 50 -17
3 U1A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 1 0
1 U
7571 0 0
2
41826.7 17
0
7 Ground~
168 86 466 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
311 0 0
2
41826.7 18
0
9 Schottky~
219 204 366 0 2 5
0 12 5
0
0 0 848 692
6 11DQ03
-22 -18 20 -10
2 D1
-8 -28 6 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
5524 0 0
2
41826.7 19
0
9 Schottky~
219 166 442 0 2 5
0 2 13
0
0 0 848 602
6 11DQ03
12 -1 54 7
2 D3
26 -11 40 -3
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
6424 0 0
2
41826.7 20
0
9 Schottky~
219 383 365 0 2 5
0 5 19
0
0 0 848 180
6 11DQ03
-22 -18 20 -10
2 D2
-8 -28 6 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
8878 0 0
2
41826.7 21
0
9 Schottky~
219 335 443 0 2 5
0 9 2
0
0 0 848 270
6 11DQ03
12 1 54 9
2 D4
26 -9 40 -1
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
3615 0 0
2
41826.7 22
0
7 Ground~
168 414 187 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7948 0 0
2
41826.7 23
0
14 Var ResistorA~
219 344 172 0 3 7
0 7 3 5
0
0 0 848 512
6 10k 1%
-22 18 20 26
2 R8
-7 8 7 16
0
0
29 %DA %1 %2 100
%DB %2 %3 9900
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
82 0 0 0 1 0 0 0
1 R
447 0 0
2
41826.7 24
0
11 Resistor:A~
219 273 71 0 2 5
0 3 4
0
0 0 880 180
3 5M1
-11 -14 10 -6
3 R15
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4827 0 0
2
41826.7 25
0
11 Resistor:A~
219 218 110 0 2 5
0 4 6
0
0 0 880 180
4 750k
-14 -14 14 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3675 0 0
2
41826.7 26
0
11 Resistor:A~
219 145 166 0 2 5
0 6 23
0
0 0 880 180
3 20k
-11 -14 10 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7278 0 0
2
41826.7 27
0
11 Resistor:A~
219 256 396 0 4 5
0 20 2 0 -1
0
0 0 880 270
3 10k
-27 2 -6 10
2 R9
-22 -10 -8 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
926 0 0
2
41826.7 28
0
11 Resistor:A~
219 208 316 0 2 5
0 18 12
0
0 0 880 180
3 10k
-10 -14 11 -6
3 R10
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6747 0 0
2
41826.7 29
0
11 Resistor:A~
219 282 316 0 2 5
0 19 18
0
0 0 880 180
3 10k
-10 -14 11 -6
3 R11
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5177 0 0
2
41826.7 30
0
11 Resistor:A~
219 335 396 0 2 5
0 19 9
0
0 0 880 270
3 10k
7 0 28 8
3 R13
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5594 0 0
2
41826.7 31
0
11 Resistor:A~
219 165 395 0 2 5
0 12 13
0
0 0 880 270
2 1k
10 0 24 8
3 R12
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9933 0 0
2
41826.7 32
0
11 Resistor:A~
219 86 396 0 4 5
0 14 2 0 -1
0
0 0 880 270
3 10k
-27 2 -6 10
2 R6
-22 -10 -8 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8987 0 0
2
41826.7 33
0
11 Resistor:A~
219 59 360 0 4 5
0 15 11 0 1
0
0 0 880 180
3 10k
-10 -14 11 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3275 0 0
2
41826.7 34
0
11 Resistor:A~
219 112 316 0 2 5
0 12 15
0
0 0 880 180
3 10k
-10 -14 11 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3551 0 0
2
41826.7 35
0
11 Resistor:A~
219 382 422 0 2 5
0 9 8
0
0 0 880 0
3 10k
-12 -14 9 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9522 0 0
2
41826.7 36
0
11 Resistor:A~
219 276 172 0 2 5
0 5 10
0
0 0 880 180
4 5.1k
-14 -14 14 -6
2 R7
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3443 0 0
2
41826.7 37
0
11 Resistor:A~
219 391 172 0 3 5
0 2 7 -1
0
0 0 880 180
4 5.1k
-14 -14 14 -6
3 R14
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3935 0 0
2
41826.7 38
0
45
1 0 3 0 0 8192 0 26 0 0 4 3
291 71
298 71
298 110
2 0 4 0 0 8320 0 26 0 0 5 3
255 71
247 71
247 110
2 0 5 0 0 8192 0 1 0 0 11 3
283 32
308 32
308 172
2 2 3 0 0 4224 0 2 25 0 0 3
286 110
346 110
346 160
1 1 4 0 0 0 0 2 27 0 0 2
268 110
236 110
1 0 6 0 0 4224 0 1 0 0 39 3
265 32
174 32
174 110
1 1 2 0 0 4096 0 24 39 0 0 3
414 181
414 172
409 172
2 1 7 0 0 4224 0 39 25 0 0 2
373 172
362 172
0 2 8 0 0 12416 0 0 37 0 0 6
244 248
4 248
4 484
416 484
416 422
400 422
1 0 9 0 0 4224 0 37 0 0 32 2
364 422
335 422
0 0 5 0 0 0 0 0 0 12 15 4
308 172
308 247
416 247
416 277
3 1 5 0 0 0 0 25 38 0 0 2
326 172
294 172
5 2 10 0 0 4224 0 5 38 0 0 2
234 172
258 172
1 2 11 0 0 4224 0 9 35 0 0 2
37 360
41 360
2 1 5 0 0 12416 0 20 22 0 0 6
216 366
244 366
244 277
416 277
416 365
392 365
2 0 12 0 0 4096 0 30 0 0 23 2
190 316
165 316
1 0 12 0 0 4096 0 20 0 0 20 2
193 366
165 366
1 1 2 0 0 0 0 15 21 0 0 2
165 460
165 452
2 2 13 0 0 4224 0 21 33 0 0 2
165 429
165 413
1 0 12 0 0 0 0 33 0 0 23 2
165 377
165 366
1 2 2 0 0 4224 0 19 34 0 0 2
86 460
86 414
1 1 14 0 0 8320 0 34 18 0 0 3
86 378
86 372
94 372
1 5 12 0 0 8320 0 36 18 0 0 4
130 316
165 316
165 366
130 366
2 0 15 0 0 8320 0 36 0 0 25 3
94 316
86 316
86 360
2 1 15 0 0 0 0 18 35 0 0 2
94 360
77 360
1 4 16 0 0 4224 0 16 18 0 0 2
112 380
112 379
1 3 17 0 0 4224 0 17 18 0 0 2
112 352
112 353
2 0 18 0 0 8320 0 12 0 0 29 3
264 359
256 359
256 316
1 2 18 0 0 0 0 30 31 0 0 2
226 316
264 316
2 0 19 0 0 4096 0 22 0 0 33 2
369 365
335 365
1 2 2 0 0 0 0 14 23 0 0 2
335 460
335 455
1 2 9 0 0 0 0 23 32 0 0 2
335 432
335 414
1 0 19 0 0 0 0 32 0 0 36 2
335 378
335 365
1 2 2 0 0 0 0 13 29 0 0 2
256 460
256 414
1 1 20 0 0 8320 0 29 12 0 0 3
256 378
256 371
264 371
1 5 19 0 0 8320 0 31 12 0 0 4
300 316
335 316
335 365
300 365
1 4 21 0 0 4224 0 10 12 0 0 2
282 379
282 378
1 3 22 0 0 4224 0 11 12 0 0 2
282 351
282 352
2 0 6 0 0 0 0 27 0 0 40 3
200 110
174 110
174 166
1 2 6 0 0 0 0 28 5 0 0 2
163 166
198 166
1 2 2 0 0 0 0 3 8 0 0 3
145 187
145 176
117 176
1 2 23 0 0 4224 0 8 28 0 0 2
117 166
127 166
1 1 2 0 0 0 0 4 5 0 0 3
190 187
190 178
198 178
1 4 24 0 0 4224 0 7 5 0 0 2
216 198
216 185
1 3 25 0 0 4224 0 6 5 0 0 2
216 145
216 159
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.25 0.001 0.001
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

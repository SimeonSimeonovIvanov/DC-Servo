CircuitMaker Text
5.6
Probes: 1
C1_2
Transient Analysis
0 369 147 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 150 10
176 83 1022 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 2 0
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 179 1190 496
9961490 0
0
6 Title:
5 Name:
0
0
0
29
10 Capacitor~
219 247 31 0 2 5
0 4 3
0
0 0 848 0
5 3.3nF
-17 -18 18 -10
2 C2
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4129 0 0
2
41825.5 0
0
7 Ground~
168 160 161 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6278 0 0
2
5.89668e-315 5.43192e-315
0
7 Ground~
168 205 161 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3482 0 0
2
5.89668e-315 5.42933e-315
0
8 Op-Amp5~
219 231 140 0 5 11
0 2 4 19 18 3
0
0 0 848 0
5 TL082
15 -25 50 -17
3 U2A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 2 0
1 U
8323 0 0
2
5.89668e-315 5.42414e-315
0
2 +V
167 231 104 0 1 3
0 19
0
0 0 53616 0
4 +15V
-14 -14 14 -6
2 V7
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3984 0 0
2
5.89668e-315 5.41896e-315
0
2 +V
167 231 181 0 1 3
0 18
0
0 0 53616 180
4 -15V
-12 -1 16 7
2 V6
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7622 0 0
2
5.89668e-315 5.41378e-315
0
11 Signal Gen~
195 101 139 0 64 64
0 17 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1120403455 -1063256064 1084227584
0 814313567 814313567 1000593163 1008981771 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 100 -5 5 0 1e-09 1e-09 0.005 0.01 0
0 0 0 0 0 0 0 0 0 0
0
0 0 1360 0
5 -5/5V
-18 -30 17 -22
2 V5
-7 -40 7 -32
8 Speed SP
-27 -40 29 -32
0
40 %D %1 %2 DC 0 PULSE(-5 5 0 1n 1n 5m 10m)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
816 0 0
2
5.89668e-315 5.4086e-315
0
7 Ground~
168 115 399 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4656 0 0
2
5.89668e-315 5.40342e-315
0
7 Ground~
168 266 397 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6356 0 0
2
5.89668e-315 5.39824e-315
0
8 Op-Amp5~
219 141 333 0 5 11
0 9 14 16 15 6
0
0 0 848 0
5 TL082
15 -25 50 -17
3 U1A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 1 0
1 U
7479 0 0
2
5.89668e-315 5.39306e-315
0
2 +V
167 141 310 0 1 3
0 16
0
0 0 53616 0
4 +15V
-14 -14 14 -6
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5690 0 0
2
5.89668e-315 5.38788e-315
0
2 +V
167 141 362 0 1 3
0 15
0
0 0 53616 180
4 -15V
-12 -1 16 7
2 V2
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5617 0 0
2
5.89668e-315 5.37752e-315
0
8 Op-Amp5~
219 297 333 0 5 11
0 10 11 12 13 7
0
0 0 848 0
5 TL082
15 -25 50 -17
3 U1B
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 5 6 8 4 7 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 2 1 0
1 U
3903 0 0
2
5.89668e-315 5.36716e-315
0
2 +V
167 297 362 0 1 3
0 13
0
0 0 53616 180
4 -15V
-12 -1 16 7
2 V3
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4452 0 0
2
5.89668e-315 5.3568e-315
0
2 +V
167 297 310 0 1 3
0 12
0
0 0 53616 0
4 +15V
-14 -14 14 -6
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6282 0 0
2
5.89668e-315 5.34643e-315
0
2 +V
167 38 329 0 1 3
0 8
0
0 0 53616 90
4 +12V
-14 -15 14 -7
2 V8
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7187 0 0
2
5.89668e-315 5.32571e-315
0
9 Schottky~
219 194 390 0 2 5
0 6 4
0
0 0 848 270
6 11DQ03
-56 2 -14 10
2 D1
-40 -10 -26 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
6866 0 0
2
5.89668e-315 5.30499e-315
0
9 Schottky~
219 349 395 0 2 5
0 4 7
0
0 0 848 90
6 11DQ03
-53 0 -11 8
2 D2
-42 -10 -28 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
7670 0 0
2
5.89668e-315 5.26354e-315
0
10 Capacitor~
219 267 74 0 2 5
0 5 3
0
0 0 848 0
4 10uF
-14 -18 14 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
951 0 0
2
5.89668e-315 0
0
11 Resistor:A~
219 219 74 0 2 5
0 5 4
0
0 0 880 180
2 1k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9536 0 0
2
5.89668e-315 5.45782e-315
0
11 Resistor:A~
219 160 134 0 2 5
0 4 17
0
0 0 880 180
2 1k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5495 0 0
2
5.89668e-315 5.45523e-315
0
11 Resistor:A~
219 141 284 0 2 5
0 6 14
0
0 0 880 180
3 10k
-10 -14 11 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8152 0 0
2
5.89668e-315 5.45264e-315
0
11 Resistor:A~
219 88 327 0 4 5
0 14 8 0 1
0
0 0 880 180
3 10k
-10 -14 11 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6223 0 0
2
5.89668e-315 5.45005e-315
0
11 Resistor:A~
219 229 366 0 2 5
0 10 3
0
0 0 880 270
3 10k
-26 2 -5 10
2 R8
-22 -10 -8 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5441 0 0
2
5.89668e-315 5.44746e-315
0
11 Resistor:A~
219 229 302 0 3 5
0 8 10 1
0
0 0 880 270
3 10k
-25 2 -4 10
2 R7
-22 -10 -8 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3189 0 0
2
5.89668e-315 5.44487e-315
0
11 Resistor:A~
219 296 284 0 2 5
0 7 11
0
0 0 880 180
3 10k
-9 -14 12 -6
3 R10
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8460 0 0
2
5.89668e-315 5.44228e-315
0
11 Resistor:A~
219 266 366 0 4 5
0 11 2 0 -1
0
0 0 880 270
3 10k
-26 2 -5 10
2 R9
-22 -10 -8 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5179 0 0
2
5.89668e-315 5.43969e-315
0
11 Resistor:A~
219 115 366 0 4 5
0 9 2 0 -1
0
0 0 880 270
3 10k
-27 2 -6 10
2 R6
-22 -10 -8 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3593 0 0
2
5.89668e-315 5.4371e-315
0
11 Resistor:A~
219 60 366 0 2 5
0 9 3
0
0 0 880 270
3 10k
-26 2 -5 10
2 R5
-22 -10 -8 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3928 0 0
2
5.89668e-315 5.43451e-315
0
35
2 0 3 0 0 4096 0 1 0 0 3 3
256 31
305 31
305 74
1 0 4 0 0 4096 0 1 0 0 5 3
238 31
189 31
189 74
2 0 3 0 0 8192 0 19 0 0 7 3
276 74
306 74
306 140
1 1 5 0 0 4224 0 19 20 0 0 2
258 74
237 74
2 0 4 0 0 8192 0 20 0 0 6 3
201 74
189 74
189 134
1 2 4 0 0 0 0 21 4 0 0 2
178 134
213 134
5 0 3 0 0 8320 0 4 0 0 16 4
249 140
370 140
370 435
229 435
0 0 4 0 0 8320 0 0 0 14 5 5
194 421
22 421
22 188
189 188
189 133
1 0 6 0 0 4224 0 17 0 0 12 2
194 379
194 330
2 0 7 0 0 4224 0 18 0 0 11 2
350 382
350 332
1 5 7 0 0 0 0 26 13 0 0 4
314 284
350 284
350 333
315 333
1 5 6 0 0 0 0 22 10 0 0 4
159 284
194 284
194 333
159 333
1 0 8 0 0 4096 0 16 0 0 15 2
49 327
61 327
2 1 4 0 0 0 0 17 18 0 0 4
194 402
194 421
350 421
350 405
2 1 8 0 0 12416 0 23 25 0 0 5
70 327
61 327
61 248
229 248
229 284
2 2 3 0 0 0 0 24 29 0 0 4
229 384
229 435
60 435
60 384
0 1 9 0 0 4224 0 0 29 20 0 3
115 339
60 339
60 348
1 2 2 0 0 4096 0 9 27 0 0 2
266 391
266 384
1 2 2 0 0 4096 0 8 28 0 0 2
115 393
115 384
1 1 9 0 0 0 0 28 10 0 0 3
115 348
115 339
123 339
1 0 10 0 0 4224 0 13 0 0 22 2
279 339
229 339
1 2 10 0 0 0 0 24 25 0 0 2
229 348
229 320
2 0 11 0 0 4096 0 13 0 0 24 2
279 327
266 327
2 1 11 0 0 8320 0 26 27 0 0 3
278 284
266 284
266 348
1 3 12 0 0 4224 0 15 13 0 0 2
297 319
297 320
1 4 13 0 0 4224 0 14 13 0 0 2
297 347
297 346
2 0 14 0 0 8320 0 22 0 0 28 3
123 284
114 284
114 327
1 2 14 0 0 0 0 23 10 0 0 2
106 327
123 327
1 4 15 0 0 4224 0 12 10 0 0 2
141 347
141 346
1 3 16 0 0 4224 0 11 10 0 0 2
141 319
141 320
1 2 2 0 0 8320 0 2 7 0 0 3
160 155
160 144
132 144
1 2 17 0 0 4224 0 7 21 0 0 2
132 134
142 134
1 1 2 0 0 0 0 3 4 0 0 3
205 155
205 146
213 146
1 4 18 0 0 4224 0 6 4 0 0 2
231 166
231 153
1 3 19 0 0 4224 0 5 4 0 0 2
231 113
231 127
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.05 0.0002 0.0002
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

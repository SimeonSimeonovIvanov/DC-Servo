CircuitMaker Text
5.6
Probes: 1
D3_A
Transient Analysis
0 263 166 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 140 10
176 83 1022 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 2 0
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 179 457 276
9961490 0
0
6 Title:
5 Name:
0
0
0
38
14 Var ResistorA~
219 301 170 0 3 7
0 20 4 5
0
0 0 832 512
7 10k 50%
-25 18 24 26
2 R1
-8 8 6 16
0
0
30 %DA %1 %2 5000
%DB %2 %3 5000
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
82 0 0 0 1 0 0 0
1 R
5130 0 0
2
41938.7 0
0
7 Ground~
168 371 185 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
391 0 0
2
41938.7 1
0
11 Signal Gen~
195 43 169 0 64 64
0 22 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1073741824 -1090519040 1056964608
0 814313567 814313567 1048576000 1056964608 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 2 -0.5 0.5 0 1e-09 1e-09 0.25 0.5 0
0 0 0 0 0 0 0 0 0 0
0
0 0 1344 0
11 -500m/500mV
-40 -30 37 -22
2 V1
-9 -40 5 -32
8 Speed SP
-27 -40 29 -32
0
49 %D %1 %2 DC 0 PULSE(-500m 500m 0 1n 1n 250m 500m)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3124 0 0
2
41938.7 2
0
2 +V
167 173 211 0 1 3
0 23
0
0 0 53600 180
4 -15V
-12 -1 16 7
2 V2
-5 -11 9 -3
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3421 0 0
2
41938.7 3
0
2 +V
167 173 134 0 1 3
0 24
0
0 0 53600 0
4 +15V
-14 -14 14 -6
2 V3
-7 -24 7 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8157 0 0
2
41938.7 4
0
8 Op-Amp5~
219 173 170 0 5 11
0 2 19 24 23 21
0
0 0 832 0
5 TL082
-39 -28 -4 -20
3 U1A
-32 -38 -11 -30
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 2 0
1 U
5572 0 0
2
41938.7 5
0
7 Ground~
168 147 191 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8901 0 0
2
41938.7 6
0
7 Ground~
168 102 191 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7361 0 0
2
41938.7 7
0
10 Capacitor~
219 234 108 0 2 5
0 3 4
0
0 0 832 0
5 220nF
-18 -18 17 -10
2 C1
-8 -28 6 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4747 0 0
2
41938.7 8
0
10 Capacitor~
219 231 30 0 2 5
0 19 5
0
0 0 832 0
5 0.1nF
-18 -18 17 -10
2 C2
-8 -28 6 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
972 0 0
2
41938.7 9
0
2 +V
167 47 299 0 1 3
0 6
0
0 0 53600 90
2 5V
-7 -15 7 -7
2 V4
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3472 0 0
2
41938.7 10
0
2 +V
167 303 331 0 1 3
0 17
0
0 0 53600 180
4 -15V
-12 -1 16 7
2 V5
-5 -11 9 -3
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9998 0 0
2
41938.7 11
0
2 +V
167 303 279 0 1 3
0 18
0
0 0 53600 0
4 +15V
-14 -14 14 -6
2 V6
-7 -24 7 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3536 0 0
2
41938.7 12
0
8 Op-Amp5~
219 303 302 0 5 11
0 16 13 18 17 14
0
0 0 832 0
5 TL082
15 -25 50 -17
3 U1B
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 5 6 8 4 7 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 2 2 0
1 U
4597 0 0
2
41938.7 13
0
7 Ground~
168 277 403 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3835 0 0
2
41938.7 14
0
7 Ground~
168 356 403 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3670 0 0
2
41938.7 15
0
7 Ground~
168 186 403 0 1 3
0 2
0
0 0 53344 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5616 0 0
2
41938.7 16
0
2 +V
167 133 332 0 1 3
0 11
0
0 0 53600 180
4 -15V
-12 -1 16 7
2 V7
-5 -11 9 -3
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9323 0 0
2
41938.7 17
0
2 +V
167 133 280 0 1 3
0 12
0
0 0 53600 0
4 +15V
-14 -14 14 -6
2 V8
-7 -24 7 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
317 0 0
2
41938.7 18
0
8 Op-Amp5~
219 133 303 0 5 11
0 9 10 12 11 7
0
0 0 832 0
5 TL082
15 -25 50 -17
3 U2A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 1 0
1 U
3108 0 0
2
41938.7 19
0
7 Ground~
168 107 403 0 1 3
0 2
0
0 0 53344 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4299 0 0
2
41938.7 20
0
9 Schottky~
219 225 303 0 2 5
0 7 5
0
0 0 832 692
6 11DQ03
-22 -18 20 -10
2 D1
-8 -28 6 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
9672 0 0
2
41938.7 21
0
9 Schottky~
219 187 379 0 2 5
0 2 8
0
0 0 832 602
6 11DQ03
12 -1 54 7
2 D2
26 -11 40 -3
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
7876 0 0
2
41938.7 22
0
9 Schottky~
219 404 302 0 2 5
0 5 14
0
0 0 832 180
6 11DQ03
-22 -18 20 -10
2 D3
-8 -28 6 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
6369 0 0
2
41938.7 23
0
9 Schottky~
219 356 380 0 2 5
0 15 2
0
0 0 832 270
6 11DQ03
12 1 54 9
2 D4
26 -9 40 -1
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
9172 0 0
2
41938.7 24
0
11 Resistor:A~
219 348 170 0 3 5
0 2 20 -1
0
0 0 864 180
4 5.1k
-14 -14 14 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7100 0 0
2
41938.7 25
0
11 Resistor:A~
219 233 170 0 2 5
0 5 21
0
0 0 864 180
4 2.7k
-14 -14 14 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3820 0 0
2
41938.7 26
0
11 Resistor:A~
219 102 164 0 2 5
0 19 22
0
0 0 864 180
3 20k
-11 -14 10 -6
2 R4
-8 -24 6 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7678 0 0
2
41938.7 27
0
11 Resistor:A~
219 175 108 0 2 5
0 3 19
0
0 0 864 180
4 220k
-14 -14 14 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
961 0 0
2
41938.7 28
0
11 Resistor:A~
219 230 69 0 2 5
0 4 3
0
0 0 864 180
3 5M1
-11 -14 10 -6
2 R6
-8 -24 6 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3178 0 0
2
41938.7 29
0
11 Resistor:A~
219 277 333 0 4 5
0 16 2 0 -1
0
0 0 864 270
4 5.1k
-30 2 -2 10
2 R7
-24 -8 -10 0
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3409 0 0
2
41938.7 30
0
11 Resistor:A~
219 229 253 0 2 5
0 13 7
0
0 0 864 180
3 10k
-10 -14 11 -6
2 R8
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3951 0 0
2
41938.7 31
0
11 Resistor:A~
219 303 253 0 2 5
0 14 13
0
0 0 864 180
3 10k
-10 -14 11 -6
2 R9
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8885 0 0
2
41938.7 32
0
11 Resistor:A~
219 356 333 0 2 5
0 14 15
0
0 0 864 270
3 10k
7 0 28 8
3 R10
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3780 0 0
2
41938.7 33
0
11 Resistor:A~
219 186 332 0 2 5
0 7 8
0
0 0 864 270
3 10k
7 0 28 8
3 R11
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9265 0 0
2
41938.7 34
0
11 Resistor:A~
219 107 333 0 4 5
0 9 2 0 -1
0
0 0 864 270
4 5.1k
-30 2 -2 10
3 R12
-27 -8 -6 0
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9442 0 0
2
41938.7 35
0
11 Resistor:A~
219 80 297 0 4 5
0 10 6 0 1
0
0 0 864 180
3 10k
-10 -14 11 -6
3 R13
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9424 0 0
2
41938.7 36
0
11 Resistor:A~
219 133 253 0 2 5
0 7 10
0
0 0 864 180
3 10k
-10 -14 11 -6
3 R14
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9968 0 0
2
41938.7 37
0
43
2 0 3 0 0 8320 0 30 0 0 30 3
212 69
204 69
204 108
1 0 4 0 0 8192 0 30 0 0 29 3
248 69
254 69
254 108
0 0 5 0 0 4096 0 0 0 34 5 2
265 170
265 216
1 2 6 0 0 4224 0 11 37 0 0 2
58 297
62 297
2 1 5 0 0 12416 0 22 24 0 0 6
237 303
265 303
265 216
437 216
437 302
413 302
2 0 7 0 0 4096 0 32 0 0 13 2
211 253
186 253
1 0 7 0 0 4096 0 22 0 0 10 2
214 303
186 303
1 1 2 0 0 4096 0 17 23 0 0 2
186 397
186 389
2 2 8 0 0 4224 0 23 35 0 0 2
186 366
186 350
1 0 7 0 0 0 0 35 0 0 13 2
186 314
186 303
1 2 2 0 0 4224 0 21 36 0 0 2
107 397
107 351
1 1 9 0 0 8320 0 36 20 0 0 3
107 315
107 309
115 309
1 5 7 0 0 8320 0 38 20 0 0 4
151 253
186 253
186 303
151 303
2 0 10 0 0 8320 0 38 0 0 15 3
115 253
107 253
107 297
2 1 10 0 0 0 0 20 37 0 0 2
115 297
98 297
1 4 11 0 0 4224 0 18 20 0 0 2
133 317
133 316
1 3 12 0 0 4224 0 19 20 0 0 2
133 289
133 290
2 0 13 0 0 8320 0 14 0 0 19 3
285 296
277 296
277 253
1 2 13 0 0 0 0 32 33 0 0 2
247 253
285 253
2 0 14 0 0 4096 0 24 0 0 23 2
390 302
356 302
1 2 2 0 0 0 0 16 25 0 0 2
356 397
356 392
1 2 15 0 0 4224 0 25 34 0 0 2
356 369
356 351
1 0 14 0 0 0 0 34 0 0 26 2
356 315
356 302
1 2 2 0 0 0 0 15 31 0 0 2
277 397
277 351
1 1 16 0 0 8320 0 31 14 0 0 3
277 315
277 308
285 308
1 5 14 0 0 8320 0 33 14 0 0 4
321 253
356 253
356 302
321 302
1 4 17 0 0 4224 0 12 14 0 0 2
303 316
303 315
1 3 18 0 0 4224 0 13 14 0 0 2
303 288
303 289
2 2 4 0 0 4224 0 9 1 0 0 3
243 108
303 108
303 158
1 1 3 0 0 0 0 9 29 0 0 2
225 108
193 108
1 0 19 0 0 4224 0 10 0 0 37 3
222 30
131 30
131 108
1 1 2 0 0 0 0 2 26 0 0 3
371 179
371 170
366 170
2 1 20 0 0 4224 0 26 1 0 0 2
330 170
319 170
2 0 5 0 0 0 0 10 0 0 35 3
240 30
265 30
265 170
3 1 5 0 0 0 0 1 27 0 0 2
283 170
251 170
5 2 21 0 0 4224 0 6 27 0 0 2
191 170
215 170
2 0 19 0 0 0 0 29 0 0 38 3
157 108
131 108
131 164
1 2 19 0 0 0 0 28 6 0 0 2
120 164
155 164
1 2 2 0 0 0 0 8 3 0 0 3
102 185
102 174
74 174
1 2 22 0 0 4224 0 3 28 0 0 2
74 164
84 164
1 1 2 0 0 0 0 7 6 0 0 3
147 185
147 176
155 176
1 4 23 0 0 4224 0 4 6 0 0 2
173 196
173 183
1 3 24 0 0 4224 0 5 6 0 0 2
173 143
173 157
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 2.5 0.01 0.01
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
